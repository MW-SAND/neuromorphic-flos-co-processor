-- ================================================================================ --
-- NEORV32 SoC - Processor-Internal Instruction Memory (IMEM)                       --
-- -------------------------------------------------------------------------------- --
-- [TIP] This file can be replaced by a technology-specific implementation to       --
--       optimize timing, area, energy, etc.                                        --
-- -------------------------------------------------------------------------------- --
-- The NEORV32 RISC-V Processor - https://github.com/stnolting/neorv32              --
-- Copyright (c) NEORV32 contributors.                                              --
-- Copyright (c) 2020 - 2024 Stephan Nolting. All rights reserved.                  --
-- Licensed under the BSD-3-Clause license, see LICENSE for details.                --
-- SPDX-License-Identifier: BSD-3-Clause                                            --
-- ================================================================================ --

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.MATH_UTILS.ALL;

library neorv32;
use neorv32.neorv32_package.all;
use neorv32.neorv32_application_image.all; -- generated by the image generator

entity neorv32_imem is
  generic (
    IMEM_SIZE    : natural; -- processor-internal instruction memory size in bytes, has to be a power of 2
    IMEM_INIT : boolean  -- implement IMEM as pre-initialized read-only memory?
  );
  port (
    clk_i     : in  std_ulogic; -- global clock line
    rstn_i    : in  std_ulogic; -- async reset, low-active
    bus_req_i : in  bus_req_t;  -- bus request
    bus_rsp_o : out bus_rsp_t   -- bus response
  );
end neorv32_imem;

architecture neorv32_imem_rtl of neorv32_imem is
  signal bus_req_i_del : bus_req_t;

  component sram is
    generic
    (
        sram_basename : string;
        banks : integer := 4;
	log2_words_per_bank : integer := 13;
        word_length : integer := 32
    );
    port 
    (
        addr : in std_logic_vector(log2(banks)+10-1 downto 0);
        din : in std_logic_vector(word_length-1 downto 0);
        we : in std_logic_vector(4-1 downto 0);
        ena : in std_logic;
        clk : in std_logic;
        dout : out std_logic_vector(word_length-1 downto 0)
    );
  end component; 

  -- alternative memory description style --
  constant alt_style_c : boolean := false; -- [TIP] enable this if synthesis fails to infer block RAM
  constant sram_c : boolean := true;

  -- local signals --
  signal rdata         : std_ulogic_vector(31 downto 0);
  signal rdata_logic   : std_logic_vector(31 downto 0);
  signal rden          : std_ulogic;
  signal addr, addr_ff : std_ulogic_vector(index_size_f(IMEM_SIZE/4)-1 downto 0);

  -- application (image) size in bytes --
  constant imem_app_size_c : natural := (application_init_image_c'length)*4;

  -- ROM - initialized with executable code --
  constant mem_rom_c : mem32_t(0 to IMEM_SIZE/4-1) := mem32_init_f(application_init_image_c, IMEM_SIZE/4);

  -- [NOTE] The memory (RAM) is built from 4 individual byte-wide memories as some synthesis tools
  --        have issues inferring 32-bit memories with individual byte-enable signals.
  -- [NOTE] Read-during-write behavior is irrelevant
  --        as read and write accesses are mutually exclusive (ensured by bus protocol).
  signal mem_ram_b0, mem_ram_b1, mem_ram_b2, mem_ram_b3 : mem8_t(0 to IMEM_SIZE/4-1);

  constant bytes_per_bank : natural := 4 * 1024; 
  constant num_banks_needed : natural := natural(index_size_f(IMEM_SIZE / bytes_per_bank)); 
  constant num_banks : natural := 2 ** num_banks_needed;

  signal sram_addr : std_logic_vector(log2(num_banks)+10-1 downto 0);
  signal sram_we : std_logic_vector(4-1 downto 0);
begin

  -- Sanity Checks --------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  assert false report
    "[NEORV32] Implementing processor-internal IMEM as " &
    cond_sel_string_f(IMEM_INIT, "pre-initialized ROM.", "blank RAM.") severity note;

  assert not ((IMEM_INIT = true) and (imem_app_size_c > IMEM_SIZE)) report
    "[NEORV32] Application image (" & natural'image(imem_app_size_c) &
    " bytes) does not fit into processor-internal IMEM (" &
    natural'image(IMEM_SIZE) & " bytes)!" severity error;


  -- Implement IMEM as pre-initialized SRAM --------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  sram_default:
  if sram_c generate
    sram_addr(index_size_f(IMEM_SIZE/4)-1 downto 0) <= std_logic_vector(addr(index_size_f(IMEM_SIZE/4)-1 downto 0));
    
    extend_sram_addr: if log2(num_banks)+10 > index_size_f(IMEM_SIZE/4) generate
      sram_addr(log2(num_banks)+10-1 downto index_size_f(IMEM_SIZE/4)) <= (others => '0');
    end generate;

    gen_write_enable: for i in 0 to 3 generate
      sram_we(i) <= bus_req_i_del.ben(i) and bus_req_i_del.rw;
    end generate;

    sram_block : sram
      generic map (
        sram_basename => "../rtl/core/hex_files/neorv32_application_image",
        banks => num_banks,
        word_length => 32,
	log2_words_per_bank => 10
      )
      port map (
        addr => sram_addr,
        din => std_logic_vector(bus_req_i_del.data),
        we => sram_we,
        ena => bus_req_i_del.stb,
        clk => clk_i,
        dout => rdata_logic
      );

    rdata <= std_ulogic_vector(rdata_logic);
    addr_ff <= (others => '0'); -- unused
  end generate;


  -- Implement IMEM as pre-initialized ROM --------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  imem_rom:
  if IMEM_INIT  and not sram_c generate

    imem_rom_default: -- default memory HDL style
    if not alt_style_c generate
      mem_access: process(clk_i)
      begin
        if rising_edge(clk_i) then
          rdata <= mem_rom_c(to_integer(unsigned(addr)));
        end if;
      end process mem_access;
      addr_ff <= (others => '0'); -- unused
    end generate;

    imem_rom_alternative: -- alternative memory HDL style
    if alt_style_c generate
      mem_access: process(clk_i)
      begin
        if rising_edge(clk_i) then
          addr_ff <= addr;
        end if;
      end process mem_access;
      rdata <= mem_rom_c(to_integer(unsigned(addr_ff)));
    end generate;

  end generate;

  -- word aligned access address --
  addr <= bus_req_i_del.addr(index_size_f(IMEM_SIZE/4)+1 downto 2);


  -- Implement IMEM as non-initialized RAM --------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  imem_ram:
  if not IMEM_INIT and not sram_c generate

    imem_ram_default: -- default memory HDL style
    if not alt_style_c generate
      mem_access: process(clk_i)
      begin
        if rising_edge(clk_i) then
          if (bus_req_i_del.stb = '1') and (bus_req_i_del.rw = '1') then
            if (bus_req_i_del.ben(0) = '1') then -- byte 0
              mem_ram_b0(to_integer(unsigned(addr))) <= bus_req_i_del.data(7 downto 0);
            end if;
            if (bus_req_i_del.ben(1) = '1') then -- byte 1
              mem_ram_b1(to_integer(unsigned(addr))) <= bus_req_i_del.data(15 downto 8);
            end if;
            if (bus_req_i_del.ben(2) = '1') then -- byte 2
              mem_ram_b2(to_integer(unsigned(addr))) <= bus_req_i_del.data(23 downto 16);
            end if;
            if (bus_req_i_del.ben(3) = '1') then -- byte 3
              mem_ram_b3(to_integer(unsigned(addr))) <= bus_req_i_del.data(31 downto 24);
            end if;
          end if;
          rdata(7  downto 0)  <= mem_ram_b0(to_integer(unsigned(addr)));
          rdata(15 downto 8)  <= mem_ram_b1(to_integer(unsigned(addr)));
          rdata(23 downto 16) <= mem_ram_b2(to_integer(unsigned(addr)));
          rdata(31 downto 24) <= mem_ram_b3(to_integer(unsigned(addr)));
        end if;
      end process mem_access;
      addr_ff <= (others => '0'); -- unused
    end generate;

    imem_ram_alternative: -- alternative memory HDL style
    if alt_style_c generate
      mem_access: process(clk_i)
      begin
        if rising_edge(clk_i) then
          addr_ff <= addr;
          if (bus_req_i_del.stb = '1') and (bus_req_i_del.rw = '1') then
            if (bus_req_i_del.ben(0) = '1') then -- byte 0
              mem_ram_b0(to_integer(unsigned(addr))) <= bus_req_i_del.data(7 downto 0);
            end if;
            if (bus_req_i_del.ben(1) = '1') then -- byte 1
              mem_ram_b1(to_integer(unsigned(addr))) <= bus_req_i_del.data(15 downto 8);
            end if;
            if (bus_req_i_del.ben(2) = '1') then -- byte 2
              mem_ram_b2(to_integer(unsigned(addr))) <= bus_req_i_del.data(23 downto 16);
            end if;
            if (bus_req_i_del.ben(3) = '1') then -- byte 3
              mem_ram_b3(to_integer(unsigned(addr))) <= bus_req_i_del.data(31 downto 24);
            end if;
          end if;
        end if;
      end process mem_access;
      rdata(7  downto 0)  <= mem_ram_b0(to_integer(unsigned(addr_ff)));
      rdata(15 downto 8)  <= mem_ram_b1(to_integer(unsigned(addr_ff)));
      rdata(23 downto 16) <= mem_ram_b2(to_integer(unsigned(addr_ff)));
      rdata(31 downto 24) <= mem_ram_b3(to_integer(unsigned(addr_ff)));
    end generate;

  end generate;


  -- Bus Response ---------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  bus_feedback: process(rstn_i, clk_i)
  begin
    if (rstn_i = '0') then
      rden          <= '0';
      bus_rsp_o.ack <= '0';
      bus_req_i_del.stb <= '0';
    elsif rising_edge(clk_i) then
      if bus_req_i_del.stb = '1' or bus_req_i.stb = '1' then
	bus_req_i_del <= bus_req_i;
      end if;

      rden <= bus_req_i_del.stb and (not bus_req_i_del.rw);
      if (IMEM_INIT = true) then
        bus_rsp_o.ack <= bus_req_i_del.stb and (not bus_req_i_del.rw); -- read-only!
      else
        bus_rsp_o.ack <= bus_req_i_del.stb;
      end if;
    end if;
  end process bus_feedback;

  bus_rsp_o.data <= rdata when (rden = '1') else (others => '0'); -- output gate
  bus_rsp_o.err  <= '0'; -- no access error possible


end neorv32_imem_rtl;
