-- Generated DMEM image with fixed point image and model weights from <MNIST_NN/model.py>
-- Image at [0x80000400, 0x8000103f]
-- Model weights at [0x80001040, 0x80008abf]
-- Built: 04.02.2025 12:13:20 (dd.mm.yyyy hh:mm:ss)
package body neorv32_dmem_image is

constant mem_ram_b0_init : mem8_t := (
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"2a",
x"5c",
x"4f",
x"4b",
x"1e",
x"12",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"6f",
x"7f",
x"7f",
x"7f",
x"7f",
x"78",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"63",
x"55",
x"1a",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"21",
x"39",
x"24",
x"39",
x"51",
x"71",
x"7f",
x"70",
x"7f",
x"7f",
x"7f",
x"7d",
x"72",
x"7f",
x"7f",
x"46",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"08",
x"21",
x"07",
x"21",
x"21",
x"21",
x"1d",
x"0a",
x"76",
x"7f",
x"35",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"29",
x"7e",
x"68",
x"09",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0b",
x"74",
x"80",
x"29",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"40",
x"7f",
x"77",
x"16",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"1d",
x"7c",
x"7f",
x"1f",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"42",
x"7f",
x"5d",
x"02",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"04",
x"66",
x"7c",
x"1d",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"3f",
x"7f",
x"5b",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"25",
x"7d",
x"78",
x"1c",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"09",
x"6e",
x"7f",
x"53",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"01",
x"65",
x"7f",
x"6d",
x"11",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"13",
x"7f",
x"7f",
x"26",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0f",
x"70",
x"7f",
x"39",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"42",
x"7f",
x"7f",
x"1a",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"1e",
x"79",
x"7f",
x"7f",
x"1a",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"3c",
x"7f",
x"7f",
x"6d",
x"14",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"3c",
x"7f",
x"67",
x"09",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"04",
x"00",
x"00",
x"02",
x"07",
x"f7",
x"ff",
x"f8",
x"05",
x"fd",
x"08",
x"fd",
x"fe",
x"00",
x"0a",
x"03",
x"0a",
x"05",
x"fc",
x"08",
x"02",
x"fb",
x"0a",
x"09",
x"ff",
x"f9",
x"f9",
x"fc",
x"f6",
x"07",
x"01",
x"fd",
x"00",
x"02",
x"01",
x"f5",
x"fb",
x"00",
x"02",
x"0a",
x"09",
x"f8",
x"01",
x"f6",
x"06",
x"f7",
x"09",
x"ff",
x"fa",
x"02",
x"00",
x"fa",
x"00",
x"ff",
x"f5",
x"07",
x"00",
x"01",
x"ff",
x"fb",
x"ff",
x"0a",
x"fb",
x"05",
x"0a",
x"f6",
x"05",
x"fd",
x"08",
x"06",
x"07",
x"fb",
x"fe",
x"fe",
x"fa",
x"f6",
x"08",
x"fd",
x"03",
x"ff",
x"fd",
x"09",
x"f9",
x"04",
x"f7",
x"f7",
x"02",
x"ff",
x"0a",
x"0a",
x"05",
x"09",
x"ff",
x"fb",
x"fc",
x"03",
x"06",
x"f9",
x"fa",
x"f6",
x"00",
x"f6",
x"09",
x"f8",
x"0a",
x"fe",
x"f8",
x"fd",
x"09",
x"ff",
x"fa",
x"03",
x"02",
x"fa",
x"f7",
x"06",
x"00",
x"fb",
x"f9",
x"08",
x"f7",
x"01",
x"e8",
x"f7",
x"f8",
x"fd",
x"0d",
x"01",
x"f7",
x"e9",
x"e8",
x"fd",
x"f8",
x"f6",
x"f6",
x"fb",
x"16",
x"f8",
x"f1",
x"f3",
x"ea",
x"04",
x"1d",
x"e9",
x"f5",
x"06",
x"e0",
x"fa",
x"ff",
x"06",
x"f8",
x"fe",
x"0c",
x"fd",
x"01",
x"f9",
x"e9",
x"fe",
x"f9",
x"07",
x"08",
x"00",
x"05",
x"02",
x"f6",
x"fc",
x"fe",
x"f9",
x"fd",
x"08",
x"03",
x"fc",
x"fd",
x"fd",
x"08",
x"03",
x"fc",
x"fe",
x"fa",
x"04",
x"fc",
x"fa",
x"02",
x"fc",
x"04",
x"09",
x"f9",
x"fc",
x"06",
x"00",
x"00",
x"05",
x"fc",
x"05",
x"09",
x"fb",
x"01",
x"08",
x"fa",
x"f9",
x"0a",
x"05",
x"ff",
x"fb",
x"00",
x"fd",
x"0a",
x"04",
x"0b",
x"0a",
x"04",
x"03",
x"09",
x"03",
x"02",
x"02",
x"ff",
x"fe",
x"06",
x"07",
x"08",
x"fe",
x"05",
x"0a",
x"fb",
x"05",
x"00",
x"0a",
x"07",
x"01",
x"f9",
x"00",
x"f6",
x"f7",
x"f8",
x"02",
x"01",
x"01",
x"fd",
x"03",
x"fd",
x"fb",
x"f7",
x"06",
x"06",
x"f8",
x"f7",
x"08",
x"fa",
x"08",
x"0a",
x"fb",
x"04",
x"ff",
x"00",
x"fb",
x"f6",
x"f8",
x"fe",
x"04",
x"fe",
x"f8",
x"08",
x"00",
x"fa",
x"ff",
x"fa",
x"06",
x"fc",
x"f6",
x"fd",
x"09",
x"f6",
x"fd",
x"fe",
x"f7",
x"ff",
x"04",
x"00",
x"f6",
x"00",
x"f8",
x"0a",
x"ff",
x"f7",
x"01",
x"03",
x"fb",
x"00",
x"fc",
x"fd",
x"fb",
x"fc",
x"fc",
x"fa",
x"07",
x"fb",
x"fe",
x"05",
x"ff",
x"f6",
x"09",
x"02",
x"07",
x"0a",
x"fb",
x"04",
x"06",
x"fd",
x"f7",
x"fb",
x"ff",
x"02",
x"01",
x"fd",
x"f6",
x"06",
x"06",
x"06",
x"03",
x"07",
x"fe",
x"eb",
x"f7",
x"fd",
x"fb",
x"0d",
x"fa",
x"01",
x"fe",
x"f7",
x"06",
x"f0",
x"fe",
x"eb",
x"03",
x"17",
x"fa",
x"00",
x"04",
x"fb",
x"02",
x"e2",
x"ec",
x"cf",
x"ec",
x"04",
x"e3",
x"fa",
x"fe",
x"f8",
x"e9",
x"e4",
x"f0",
x"c2",
x"00",
x"17",
x"ec",
x"02",
x"fa",
x"01",
x"e8",
x"f0",
x"f5",
x"d2",
x"01",
x"21",
x"f3",
x"ec",
x"ee",
x"dc",
x"e8",
x"eb",
x"e4",
x"d2",
x"ed",
x"10",
x"e6",
x"e4",
x"e6",
x"d1",
x"ec",
x"d3",
x"f6",
x"c8",
x"e7",
x"0d",
x"e3",
x"e9",
x"eb",
x"22",
x"ee",
x"d1",
x"eb",
x"ae",
x"ee",
x"08",
x"dd",
x"cf",
x"df",
x"1a",
x"ee",
x"c0",
x"e4",
x"b3",
x"d7",
x"1b",
x"d6",
x"be",
x"c2",
x"23",
x"d3",
x"bd",
x"e7",
x"c3",
x"e0",
x"22",
x"d6",
x"cd",
x"cc",
x"d7",
x"0c",
x"e5",
x"dc",
x"df",
x"cf",
x"e9",
x"dd",
x"cc",
x"da",
x"15",
x"12",
x"fb",
x"e3",
x"b7",
x"c5",
x"f3",
x"d2",
x"d9",
x"d8",
x"0f",
x"d6",
x"16",
x"ca",
x"b5",
x"c8",
x"ea",
x"dd",
x"db",
x"d7",
x"1b",
x"c4",
x"ee",
x"cd",
x"a6",
x"be",
x"10",
x"e3",
x"d9",
x"c0",
x"ec",
x"e8",
x"c8",
x"e0",
x"c0",
x"cd",
x"5c",
x"f3",
x"dd",
x"e3",
x"e3",
x"01",
x"b8",
x"e4",
x"bf",
x"c6",
x"3b",
x"fe",
x"d7",
x"d5",
x"ef",
x"03",
x"cc",
x"dd",
x"c5",
x"d1",
x"27",
x"04",
x"d8",
x"d8",
x"f4",
x"fc",
x"de",
x"e9",
x"d8",
x"e8",
x"1d",
x"f9",
x"e9",
x"eb",
x"02",
x"f3",
x"dd",
x"f3",
x"e1",
x"df",
x"19",
x"f3",
x"f4",
x"ea",
x"fc",
x"05",
x"e9",
x"05",
x"de",
x"f6",
x"1a",
x"f6",
x"f4",
x"e1",
x"0b",
x"f9",
x"06",
x"09",
x"f6",
x"fd",
x"03",
x"03",
x"fd",
x"f8",
x"f9",
x"0a",
x"03",
x"fb",
x"00",
x"04",
x"f6",
x"fb",
x"00",
x"06",
x"06",
x"f8",
x"ff",
x"02",
x"f5",
x"fc",
x"fa",
x"fc",
x"f9",
x"00",
x"f6",
x"08",
x"09",
x"fd",
x"0a",
x"04",
x"f7",
x"fe",
x"f7",
x"fc",
x"0a",
x"fe",
x"04",
x"01",
x"09",
x"04",
x"00",
x"fb",
x"fb",
x"00",
x"fb",
x"09",
x"05",
x"06",
x"fa",
x"f8",
x"01",
x"00",
x"02",
x"ff",
x"07",
x"fb",
x"05",
x"00",
x"f9",
x"01",
x"16",
x"04",
x"f3",
x"fc",
x"19",
x"fe",
x"e2",
x"ef",
x"e2",
x"e5",
x"03",
x"f2",
x"f2",
x"ef",
x"12",
x"00",
x"e9",
x"f9",
x"e3",
x"e6",
x"1b",
x"ef",
x"f8",
x"e1",
x"f4",
x"e7",
x"eb",
x"e4",
x"e4",
x"f0",
x"08",
x"f4",
x"f5",
x"fc",
x"e6",
x"e6",
x"e7",
x"ef",
x"c8",
x"ec",
x"17",
x"ed",
x"e5",
x"e9",
x"e4",
x"e1",
x"df",
x"d7",
x"b7",
x"eb",
x"2b",
x"db",
x"d2",
x"e0",
x"bf",
x"d5",
x"f2",
x"c4",
x"9e",
x"e0",
x"17",
x"e7",
x"c3",
x"f2",
x"cc",
x"db",
x"fb",
x"af",
x"9d",
x"c2",
x"16",
x"e2",
x"9b",
x"dd",
x"cb",
x"c4",
x"e0",
x"e0",
x"87",
x"bc",
x"27",
x"d4",
x"96",
x"cd",
x"b4",
x"ce",
x"e8",
x"fd",
x"5f",
x"c7",
x"20",
x"cc",
x"6f",
x"bc",
x"bd",
x"f4",
x"f8",
x"fc",
x"87",
x"9c",
x"21",
x"cc",
x"85",
x"b1",
x"b2",
x"27",
x"e9",
x"f1",
x"b5",
x"71",
x"19",
x"c1",
x"64",
x"95",
x"90",
x"1f",
x"d7",
x"05",
x"bb",
x"66",
x"0a",
x"d2",
x"59",
x"9d",
x"75",
x"29",
x"e4",
x"d8",
x"9f",
x"b7",
x"07",
x"c8",
x"51",
x"a7",
x"aa",
x"1f",
x"e6",
x"ee",
x"9e",
x"d8",
x"16",
x"ce",
x"43",
x"a7",
x"95",
x"f7",
x"dc",
x"e9",
x"b5",
x"dd",
x"1c",
x"e5",
x"98",
x"ab",
x"96",
x"f0",
x"d3",
x"d8",
x"62",
x"e0",
x"1d",
x"ea",
x"d6",
x"98",
x"b0",
x"02",
x"c1",
x"bd",
x"9c",
x"e0",
x"1f",
x"e6",
x"64",
x"af",
x"97",
x"f8",
x"b6",
x"a9",
x"ac",
x"d2",
x"2e",
x"fb",
x"81",
x"cc",
x"b5",
x"e5",
x"d0",
x"cc",
x"bf",
x"cd",
x"3a",
x"fd",
x"92",
x"d9",
x"bb",
x"d8",
x"ad",
x"d8",
x"cd",
x"e6",
x"3e",
x"ec",
x"a7",
x"ec",
x"d7",
x"e4",
x"f1",
x"d9",
x"c4",
x"d8",
x"38",
x"e6",
x"d9",
x"e4",
x"eb",
x"f1",
x"26",
x"ee",
x"dc",
x"ca",
x"fa",
x"f3",
x"d9",
x"e9",
x"e6",
x"fb",
x"1f",
x"f6",
x"e8",
x"d9",
x"ed",
x"06",
x"ee",
x"ff",
x"06",
x"00",
x"00",
x"fc",
x"00",
x"02",
x"f9",
x"0a",
x"04",
x"fb",
x"fb",
x"09",
x"06",
x"05",
x"f9",
x"03",
x"fc",
x"fa",
x"09",
x"06",
x"00",
x"0b",
x"02",
x"ff",
x"fc",
x"07",
x"09",
x"f6",
x"fe",
x"f7",
x"fd",
x"0a",
x"f7",
x"fd",
x"fe",
x"00",
x"f6",
x"fd",
x"07",
x"fb",
x"ff",
x"1d",
x"ed",
x"e6",
x"f7",
x"ea",
x"e6",
x"f7",
x"eb",
x"06",
x"01",
x"23",
x"e8",
x"ec",
x"e0",
x"00",
x"0e",
x"e3",
x"e8",
x"de",
x"f1",
x"e5",
x"ce",
x"dd",
x"d1",
x"1b",
x"28",
x"e0",
x"e5",
x"e9",
x"f0",
x"d8",
x"05",
x"23",
x"dd",
x"cf",
x"18",
x"dc",
x"cf",
x"dc",
x"c6",
x"e3",
x"fc",
x"fb",
x"be",
x"b7",
x"1d",
x"df",
x"c9",
x"dd",
x"bc",
x"e7",
x"0a",
x"01",
x"cd",
x"c5",
x"0e",
x"b6",
x"9c",
x"d6",
x"f0",
x"ba",
x"00",
x"06",
x"b3",
x"d1",
x"01",
x"c8",
x"de",
x"ca",
x"c4",
x"d8",
x"2a",
x"e5",
x"9c",
x"e1",
x"09",
x"b8",
x"d8",
x"c2",
x"c0",
x"b6",
x"10",
x"f0",
x"9f",
x"e8",
x"04",
x"c5",
x"e2",
x"a3",
x"d8",
x"ae",
x"09",
x"ff",
x"ae",
x"cf",
x"f6",
x"a3",
x"c7",
x"a6",
x"cf",
x"d5",
x"fc",
x"0e",
x"83",
x"f3",
x"f5",
x"ba",
x"c1",
x"89",
x"f8",
x"d9",
x"19",
x"ff",
x"6d",
x"f3",
x"f9",
x"a6",
x"d4",
x"6f",
x"ea",
x"d2",
x"fe",
x"07",
x"a6",
x"ef",
x"03",
x"be",
x"c3",
x"61",
x"ec",
x"f0",
x"fc",
x"11",
x"ab",
x"f3",
x"ff",
x"bf",
x"cf",
x"65",
x"ea",
x"fb",
x"00",
x"fe",
x"c0",
x"dd",
x"f9",
x"c5",
x"bf",
x"76",
x"e8",
x"f0",
x"f8",
x"10",
x"c4",
x"ef",
x"00",
x"c4",
x"bc",
x"93",
x"d2",
x"ce",
x"ea",
x"0c",
x"b8",
x"f6",
x"ff",
x"e2",
x"d0",
x"cf",
x"d4",
x"ee",
x"f0",
x"13",
x"dd",
x"ec",
x"19",
x"dc",
x"c1",
x"a3",
x"e7",
x"d8",
x"e8",
x"31",
x"ea",
x"04",
x"fb",
x"e9",
x"db",
x"a6",
x"cc",
x"e3",
x"fa",
x"06",
x"e0",
x"fe",
x"09",
x"e0",
x"ef",
x"c9",
x"ce",
x"da",
x"f0",
x"c1",
x"ee",
x"fd",
x"0d",
x"e5",
x"00",
x"dd",
x"e4",
x"bb",
x"a5",
x"b4",
x"de",
x"d5",
x"0b",
x"ef",
x"1e",
x"de",
x"ea",
x"aa",
x"0e",
x"c6",
x"c1",
x"ea",
x"22",
x"ea",
x"fe",
x"ee",
x"f2",
x"ca",
x"1e",
x"fa",
x"f4",
x"ff",
x"e7",
x"f6",
x"f5",
x"f2",
x"f1",
x"d3",
x"e9",
x"f8",
x"e9",
x"fe",
x"16",
x"fb",
x"e7",
x"f6",
x"05",
x"02",
x"06",
x"03",
x"08",
x"f8",
x"fa",
x"f6",
x"04",
x"fc",
x"03",
x"f7",
x"fd",
x"06",
x"08",
x"04",
x"02",
x"00",
x"06",
x"00",
x"00",
x"fa",
x"f1",
x"1c",
x"f6",
x"f4",
x"fb",
x"01",
x"f4",
x"fc",
x"fe",
x"15",
x"d4",
x"f7",
x"e8",
x"e8",
x"e1",
x"02",
x"04",
x"f2",
x"e3",
x"f8",
x"d8",
x"18",
x"d4",
x"ee",
x"e9",
x"0e",
x"d2",
x"e7",
x"c6",
x"09",
x"cd",
x"0f",
x"02",
x"ad",
x"13",
x"f9",
x"d3",
x"e6",
x"ac",
x"12",
x"f7",
x"30",
x"f0",
x"af",
x"07",
x"d0",
x"b6",
x"db",
x"c5",
x"f7",
x"1c",
x"11",
x"d9",
x"e0",
x"e8",
x"aa",
x"b9",
x"c9",
x"e7",
x"fc",
x"05",
x"02",
x"e9",
x"e4",
x"f8",
x"a3",
x"f2",
x"d4",
x"f9",
x"fa",
x"00",
x"0d",
x"cb",
x"d7",
x"00",
x"9d",
x"fc",
x"ae",
x"01",
x"e9",
x"1b",
x"12",
x"dd",
x"e5",
x"ec",
x"99",
x"00",
x"87",
x"fa",
x"ea",
x"0c",
x"0b",
x"cf",
x"f7",
x"fc",
x"7b",
x"06",
x"bf",
x"f5",
x"df",
x"ff",
x"08",
x"d9",
x"05",
x"e2",
x"c7",
x"f5",
x"cd",
x"f3",
x"e9",
x"11",
x"0d",
x"e8",
x"f3",
x"e1",
x"cf",
x"fa",
x"c9",
x"f8",
x"00",
x"02",
x"09",
x"e8",
x"e3",
x"e3",
x"d2",
x"fd",
x"c4",
x"ee",
x"f8",
x"12",
x"01",
x"e1",
x"f6",
x"e9",
x"c9",
x"fe",
x"c3",
x"fd",
x"f1",
x"fc",
x"0a",
x"ce",
x"0a",
x"e8",
x"a5",
x"ff",
x"be",
x"eb",
x"f6",
x"05",
x"04",
x"e8",
x"05",
x"ec",
x"87",
x"fe",
x"ac",
x"fd",
x"ee",
x"f6",
x"ee",
x"e7",
x"f6",
x"01",
x"4b",
x"ea",
x"b1",
x"fe",
x"e5",
x"f0",
x"0b",
x"d8",
x"03",
x"f2",
x"69",
x"f8",
x"ba",
x"f6",
x"08",
x"ec",
x"fd",
x"ff",
x"ff",
x"fb",
x"6f",
x"f8",
x"a3",
x"f9",
x"ff",
x"ec",
x"f4",
x"0c",
x"ea",
x"01",
x"79",
x"f5",
x"bc",
x"e4",
x"fa",
x"d8",
x"eb",
x"14",
x"0c",
x"03",
x"ec",
x"fb",
x"5b",
x"f5",
x"ee",
x"c7",
x"fd",
x"1b",
x"01",
x"10",
x"db",
x"ed",
x"93",
x"fa",
x"ec",
x"b2",
x"97",
x"17",
x"16",
x"04",
x"d0",
x"e4",
x"a4",
x"d6",
x"b6",
x"ce",
x"a6",
x"26",
x"1c",
x"fe",
x"e2",
x"0c",
x"cd",
x"d8",
x"a3",
x"02",
x"d8",
x"04",
x"07",
x"ed",
x"f6",
x"19",
x"dc",
x"d5",
x"d0",
x"dd",
x"f1",
x"e5",
x"f9",
x"0f",
x"f6",
x"0b",
x"ed",
x"f3",
x"e4",
x"e9",
x"fb",
x"dd",
x"cb",
x"19",
x"ef",
x"02",
x"e8",
x"04",
x"fa",
x"0a",
x"f6",
x"01",
x"fa",
x"04",
x"fe",
x"f7",
x"fe",
x"f6",
x"f9",
x"f9",
x"fb",
x"04",
x"02",
x"fa",
x"fa",
x"f8",
x"07",
x"da",
x"09",
x"ee",
x"eb",
x"ce",
x"cc",
x"0a",
x"e6",
x"df",
x"de",
x"da",
x"1d",
x"ec",
x"19",
x"f4",
x"f0",
x"c9",
x"11",
x"d1",
x"dd",
x"ca",
x"2c",
x"fb",
x"16",
x"00",
x"9e",
x"06",
x"d0",
x"bf",
x"de",
x"c3",
x"1b",
x"03",
x"16",
x"03",
x"cc",
x"f7",
x"0d",
x"cb",
x"ce",
x"00",
x"15",
x"f6",
x"0e",
x"fa",
x"dd",
x"e0",
x"01",
x"f0",
x"ad",
x"fb",
x"f5",
x"f7",
x"13",
x"f2",
x"f5",
x"e9",
x"05",
x"f6",
x"a3",
x"fb",
x"d6",
x"01",
x"05",
x"f6",
x"ed",
x"05",
x"fc",
x"ee",
x"c7",
x"f7",
x"d2",
x"fc",
x"03",
x"ff",
x"fe",
x"e7",
x"05",
x"f1",
x"cf",
x"05",
x"e8",
x"04",
x"08",
x"f9",
x"ff",
x"ff",
x"fe",
x"ed",
x"df",
x"05",
x"d5",
x"0e",
x"ff",
x"f5",
x"f9",
x"de",
x"f1",
x"02",
x"09",
x"ef",
x"d4",
x"01",
x"09",
x"f4",
x"f8",
x"f0",
x"f8",
x"08",
x"04",
x"10",
x"f0",
x"0c",
x"00",
x"e9",
x"f8",
x"e9",
x"ff",
x"fd",
x"fc",
x"09",
x"f0",
x"03",
x"ff",
x"f9",
x"f5",
x"f2",
x"fa",
x"0b",
x"f0",
x"06",
x"fb",
x"0c",
x"02",
x"0b",
x"f0",
x"e7",
x"e5",
x"05",
x"ea",
x"04",
x"e9",
x"0d",
x"04",
x"14",
x"fc",
x"f1",
x"e8",
x"03",
x"d0",
x"02",
x"e1",
x"0a",
x"f4",
x"07",
x"01",
x"ed",
x"c6",
x"0f",
x"d9",
x"0b",
x"f3",
x"09",
x"f5",
x"10",
x"0c",
x"0b",
x"ca",
x"00",
x"d6",
x"fd",
x"f3",
x"fc",
x"fd",
x"04",
x"f8",
x"0d",
x"b2",
x"fd",
x"da",
x"f8",
x"fa",
x"f4",
x"f7",
x"00",
x"0c",
x"0f",
x"90",
x"f8",
x"d9",
x"f8",
x"10",
x"04",
x"ee",
x"fe",
x"09",
x"00",
x"b3",
x"f7",
x"cb",
x"f9",
x"1a",
x"04",
x"ee",
x"0c",
x"14",
x"f6",
x"bb",
x"f4",
x"98",
x"f3",
x"0f",
x"de",
x"d4",
x"0e",
x"0b",
x"0a",
x"7d",
x"e0",
x"56",
x"d0",
x"fe",
x"bc",
x"ca",
x"f4",
x"19",
x"fb",
x"ac",
x"e5",
x"72",
x"a9",
x"a6",
x"fc",
x"b3",
x"da",
x"18",
x"ea",
x"da",
x"01",
x"ad",
x"ae",
x"cf",
x"d1",
x"e4",
x"cf",
x"15",
x"0b",
x"de",
x"f6",
x"d9",
x"f1",
x"eb",
x"e2",
x"e9",
x"da",
x"f4",
x"20",
x"ee",
x"f1",
x"ee",
x"07",
x"04",
x"fc",
x"01",
x"fd",
x"01",
x"01",
x"06",
x"fd",
x"fe",
x"fd",
x"03",
x"f2",
x"1b",
x"08",
x"f7",
x"09",
x"02",
x"eb",
x"eb",
x"e2",
x"d8",
x"fa",
x"f2",
x"d3",
x"19",
x"f1",
x"29",
x"cd",
x"d7",
x"da",
x"12",
x"ee",
x"28",
x"d1",
x"a5",
x"ac",
x"20",
x"cb",
x"cb",
x"ca",
x"20",
x"00",
x"07",
x"0b",
x"da",
x"ff",
x"01",
x"cd",
x"af",
x"03",
x"f9",
x"09",
x"09",
x"07",
x"fa",
x"00",
x"f6",
x"fe",
x"88",
x"01",
x"fa",
x"00",
x"14",
x"fe",
x"fa",
x"e9",
x"15",
x"f3",
x"cf",
x"f5",
x"e6",
x"0a",
x"fe",
x"05",
x"f5",
x"fa",
x"10",
x"f2",
x"ca",
x"f2",
x"db",
x"04",
x"02",
x"fd",
x"f4",
x"fc",
x"11",
x"f5",
x"e8",
x"cf",
x"d4",
x"08",
x"0b",
x"fc",
x"f4",
x"f0",
x"09",
x"fb",
x"f2",
x"fd",
x"e3",
x"ff",
x"0f",
x"e8",
x"fe",
x"df",
x"13",
x"ec",
x"f3",
x"f0",
x"f6",
x"03",
x"03",
x"e1",
x"02",
x"f8",
x"1b",
x"fe",
x"09",
x"fa",
x"f2",
x"00",
x"0a",
x"e3",
x"ff",
x"ee",
x"13",
x"05",
x"0b",
x"0e",
x"e9",
x"05",
x"0b",
x"d9",
x"00",
x"eb",
x"f9",
x"03",
x"24",
x"02",
x"f0",
x"00",
x"01",
x"dc",
x"00",
x"e9",
x"f9",
x"fb",
x"1a",
x"fc",
x"de",
x"06",
x"08",
x"d2",
x"f7",
x"f5",
x"f5",
x"0d",
x"14",
x"07",
x"df",
x"09",
x"08",
x"d6",
x"f4",
x"e2",
x"0b",
x"03",
x"20",
x"06",
x"e1",
x"fe",
x"00",
x"e0",
x"fb",
x"f7",
x"08",
x"01",
x"16",
x"0c",
x"f7",
x"fe",
x"0a",
x"e1",
x"f8",
x"e5",
x"f6",
x"f7",
x"15",
x"05",
x"f2",
x"f3",
x"ee",
x"ec",
x"0a",
x"f2",
x"fd",
x"01",
x"04",
x"02",
x"f9",
x"ee",
x"04",
x"f9",
x"0c",
x"f1",
x"f4",
x"00",
x"06",
x"07",
x"fd",
x"fb",
x"ff",
x"f6",
x"fc",
x"f8",
x"0c",
x"00",
x"f3",
x"19",
x"f9",
x"f7",
x"f2",
x"0a",
x"0d",
x"fe",
x"fc",
x"f6",
x"df",
x"ec",
x"03",
x"d9",
x"e7",
x"25",
x"0f",
x"fa",
x"c8",
x"01",
x"ca",
x"b3",
x"ee",
x"bd",
x"e1",
x"f8",
x"30",
x"e4",
x"cf",
x"e3",
x"ad",
x"6b",
x"7e",
x"d8",
x"97",
x"d5",
x"20",
x"f6",
x"a8",
x"01",
x"cf",
x"a8",
x"c8",
x"e2",
x"cb",
x"08",
x"1a",
x"e1",
x"ac",
x"fe",
x"bf",
x"e0",
x"e7",
x"e5",
x"f8",
x"db",
x"02",
x"13",
x"d5",
x"e8",
x"e6",
x"06",
x"08",
x"ee",
x"fd",
x"02",
x"f7",
x"01",
x"01",
x"06",
x"f4",
x"d4",
x"d5",
x"cf",
x"39",
x"eb",
x"e2",
x"f3",
x"18",
x"ce",
x"c3",
x"e4",
x"e2",
x"19",
x"d1",
x"cc",
x"fe",
x"eb",
x"28",
x"c1",
x"d4",
x"e1",
x"d0",
x"05",
x"0d",
x"ee",
x"a2",
x"b4",
x"26",
x"b0",
x"d0",
x"ba",
x"06",
x"0a",
x"16",
x"09",
x"a5",
x"f1",
x"ef",
x"f2",
x"92",
x"f9",
x"d2",
x"01",
x"0e",
x"1f",
x"df",
x"f9",
x"fa",
x"eb",
x"b4",
x"fb",
x"cb",
x"06",
x"03",
x"00",
x"f2",
x"e9",
x"07",
x"f0",
x"d4",
x"00",
x"f5",
x"fc",
x"fe",
x"01",
x"00",
x"fd",
x"1b",
x"00",
x"d5",
x"d8",
x"da",
x"0a",
x"00",
x"fd",
x"01",
x"fb",
x"0a",
x"07",
x"f1",
x"ff",
x"e4",
x"fb",
x"00",
x"00",
x"fd",
x"f9",
x"0d",
x"01",
x"f6",
x"fa",
x"f5",
x"fb",
x"fb",
x"f7",
x"05",
x"f5",
x"1c",
x"05",
x"fa",
x"04",
x"e9",
x"07",
x"01",
x"fb",
x"07",
x"f5",
x"0d",
x"f8",
x"01",
x"f7",
x"f6",
x"fd",
x"06",
x"e1",
x"07",
x"f1",
x"11",
x"ff",
x"14",
x"08",
x"f3",
x"08",
x"06",
x"e2",
x"f5",
x"e5",
x"0b",
x"f3",
x"1e",
x"0a",
x"ee",
x"00",
x"0e",
x"d4",
x"02",
x"f8",
x"f7",
x"f4",
x"24",
x"03",
x"e5",
x"00",
x"0a",
x"d7",
x"ec",
x"f6",
x"f6",
x"0b",
x"33",
x"01",
x"ef",
x"fd",
x"00",
x"d6",
x"fa",
x"e7",
x"09",
x"ff",
x"23",
x"14",
x"ed",
x"ea",
x"08",
x"e9",
x"01",
x"e6",
x"0b",
x"f3",
x"12",
x"14",
x"ef",
x"f4",
x"f8",
x"f4",
x"00",
x"de",
x"13",
x"00",
x"01",
x"0f",
x"fa",
x"fa",
x"08",
x"fa",
x"fd",
x"dc",
x"08",
x"fb",
x"fc",
x"02",
x"02",
x"fd",
x"fd",
x"f6",
x"00",
x"e2",
x"12",
x"04",
x"03",
x"fc",
x"00",
x"ff",
x"ef",
x"03",
x"0e",
x"e3",
x"13",
x"0b",
x"00",
x"fe",
x"00",
x"1a",
x"ee",
x"0b",
x"04",
x"e3",
x"11",
x"01",
x"e9",
x"02",
x"f7",
x"c9",
x"ea",
x"0f",
x"1b",
x"d7",
x"07",
x"0e",
x"ec",
x"ca",
x"c6",
x"aa",
x"ac",
x"f7",
x"30",
x"ff",
x"f1",
x"f6",
x"c0",
x"9e",
x"82",
x"e3",
x"93",
x"f0",
x"3f",
x"ed",
x"c5",
x"dd",
x"c0",
x"a2",
x"dd",
x"e4",
x"d4",
x"0a",
x"00",
x"05",
x"b0",
x"ef",
x"9a",
x"d2",
x"f1",
x"eb",
x"f7",
x"cb",
x"08",
x"02",
x"e4",
x"f3",
x"d3",
x"24",
x"04",
x"dd",
x"f2",
x"d3",
x"f7",
x"fe",
x"e9",
x"f5",
x"eb",
x"d4",
x"d2",
x"00",
x"e7",
x"cf",
x"d9",
x"03",
x"41",
x"c9",
x"d9",
x"09",
x"e8",
x"05",
x"af",
x"f4",
x"c7",
x"e4",
x"20",
x"9f",
x"c2",
x"fe",
x"d6",
x"f5",
x"01",
x"f9",
x"97",
x"93",
x"24",
x"f2",
x"a8",
x"c4",
x"f8",
x"11",
x"16",
x"fb",
x"a2",
x"f3",
x"fd",
x"f4",
x"d8",
x"ef",
x"ca",
x"fb",
x"0f",
x"13",
x"e7",
x"f0",
x"09",
x"fa",
x"e5",
x"00",
x"cd",
x"fd",
x"fe",
x"00",
x"f1",
x"e4",
x"0a",
x"04",
x"ec",
x"f8",
x"f2",
x"f6",
x"fc",
x"ff",
x"f0",
x"f0",
x"26",
x"0e",
x"e5",
x"fb",
x"dd",
x"02",
x"02",
x"f1",
x"07",
x"fa",
x"16",
x"01",
x"ff",
x"0f",
x"dd",
x"fc",
x"f8",
x"fb",
x"00",
x"f3",
x"0b",
x"0b",
x"f1",
x"fb",
x"f0",
x"10",
x"00",
x"f2",
x"0a",
x"f0",
x"0e",
x"03",
x"f3",
x"f5",
x"f1",
x"0a",
x"00",
x"f6",
x"04",
x"fd",
x"1e",
x"ff",
x"ec",
x"0b",
x"f8",
x"fd",
x"0b",
x"ea",
x"00",
x"ed",
x"12",
x"04",
x"f3",
x"fe",
x"01",
x"fb",
x"fd",
x"e7",
x"f5",
x"f6",
x"02",
x"0a",
x"05",
x"02",
x"00",
x"05",
x"03",
x"d7",
x"f2",
x"e0",
x"06",
x"f4",
x"18",
x"15",
x"f5",
x"fa",
x"02",
x"dc",
x"eb",
x"db",
x"15",
x"f5",
x"14",
x"1d",
x"e8",
x"f6",
x"04",
x"ea",
x"f6",
x"db",
x"0f",
x"00",
x"0a",
x"19",
x"01",
x"00",
x"00",
x"f1",
x"fe",
x"de",
x"11",
x"f5",
x"04",
x"10",
x"f9",
x"f2",
x"12",
x"fa",
x"f6",
x"ca",
x"12",
x"ff",
x"fb",
x"0b",
x"f9",
x"06",
x"0a",
x"fc",
x"09",
x"c5",
x"01",
x"08",
x"f7",
x"02",
x"eb",
x"04",
x"0b",
x"fb",
x"13",
x"cd",
x"0e",
x"02",
x"f6",
x"10",
x"e7",
x"f6",
x"04",
x"fc",
x"13",
x"d7",
x"f6",
x"06",
x"0b",
x"fa",
x"e9",
x"02",
x"09",
x"fa",
x"03",
x"d0",
x"0c",
x"11",
x"fa",
x"05",
x"d9",
x"07",
x"c7",
x"04",
x"18",
x"ad",
x"0f",
x"0d",
x"e8",
x"db",
x"9b",
x"80",
x"73",
x"ec",
x"42",
x"aa",
x"e8",
x"00",
x"e1",
x"75",
x"84",
x"6f",
x"80",
x"f0",
x"40",
x"bc",
x"b9",
x"e3",
x"d7",
x"95",
x"d6",
x"de",
x"c6",
x"eb",
x"09",
x"fa",
x"9d",
x"0a",
x"8c",
x"e4",
x"ee",
x"f1",
x"ee",
x"e5",
x"f7",
x"de",
x"e3",
x"26",
x"dd",
x"f4",
x"ef",
x"f6",
x"e9",
x"fb",
x"00",
x"01",
x"0d",
x"f1",
x"f1",
x"ed",
x"e2",
x"dc",
x"df",
x"d4",
x"ef",
x"fa",
x"24",
x"c8",
x"d1",
x"05",
x"e0",
x"e3",
x"db",
x"fe",
x"d2",
x"d1",
x"1d",
x"b2",
x"c4",
x"f2",
x"d2",
x"00",
x"05",
x"d6",
x"96",
x"a8",
x"1f",
x"e2",
x"ca",
x"e1",
x"eb",
x"fd",
x"1c",
x"e9",
x"c3",
x"08",
x"1a",
x"e3",
x"c1",
x"f6",
x"ba",
x"13",
x"fd",
x"f9",
x"e3",
x"df",
x"0b",
x"0d",
x"ee",
x"f8",
x"e9",
x"fa",
x"0c",
x"ef",
x"ff",
x"fc",
x"0f",
x"0b",
x"06",
x"f9",
x"08",
x"05",
x"0d",
x"03",
x"fd",
x"07",
x"0a",
x"0e",
x"f6",
x"f8",
x"00",
x"f4",
x"fa",
x"fb",
x"0f",
x"ff",
x"0c",
x"0b",
x"f9",
x"ff",
x"e1",
x"0b",
x"f7",
x"fa",
x"02",
x"f0",
x"05",
x"0a",
x"f6",
x"04",
x"fd",
x"03",
x"ee",
x"ed",
x"06",
x"eb",
x"ff",
x"05",
x"01",
x"fa",
x"03",
x"02",
x"e2",
x"f4",
x"1e",
x"fa",
x"0c",
x"0c",
x"00",
x"02",
x"01",
x"05",
x"e3",
x"ec",
x"08",
x"f5",
x"1f",
x"03",
x"f9",
x"13",
x"fd",
x"00",
x"f8",
x"f4",
x"fd",
x"e6",
x"0c",
x"ff",
x"01",
x"00",
x"17",
x"05",
x"0b",
x"d8",
x"ed",
x"f0",
x"19",
x"ef",
x"0e",
x"00",
x"21",
x"0a",
x"10",
x"de",
x"e5",
x"d8",
x"13",
x"e1",
x"06",
x"19",
x"0f",
x"07",
x"16",
x"fa",
x"e3",
x"de",
x"0c",
x"f9",
x"fb",
x"19",
x"fd",
x"05",
x"08",
x"f7",
x"e9",
x"c4",
x"1e",
x"02",
x"f0",
x"14",
x"02",
x"03",
x"08",
x"fa",
x"f7",
x"cd",
x"0a",
x"f7",
x"f7",
x"12",
x"e6",
x"00",
x"05",
x"f9",
x"e7",
x"d6",
x"12",
x"05",
x"f4",
x"09",
x"e8",
x"f5",
x"16",
x"00",
x"f7",
x"e8",
x"02",
x"00",
x"ff",
x"00",
x"f6",
x"f3",
x"10",
x"00",
x"17",
x"e1",
x"07",
x"13",
x"f0",
x"00",
x"ed",
x"06",
x"20",
x"f7",
x"12",
x"e1",
x"12",
x"11",
x"ee",
x"19",
x"ce",
x"09",
x"ea",
x"fe",
x"28",
x"ec",
x"03",
x"16",
x"e7",
x"e2",
x"b9",
x"87",
x"22",
x"d1",
x"58",
x"cf",
x"e7",
x"f6",
x"d4",
x"8b",
x"a4",
x"92",
x"ba",
x"d6",
x"66",
x"9b",
x"e7",
x"ee",
x"ca",
x"8b",
x"de",
x"e7",
x"d7",
x"d3",
x"22",
x"c2",
x"fc",
x"1d",
x"9a",
x"df",
x"ee",
x"de",
x"ee",
x"d2",
x"0e",
x"d7",
x"1a",
x"d9",
x"dd",
x"fe",
x"00",
x"f1",
x"f6",
x"ee",
x"ee",
x"f8",
x"17",
x"ec",
x"e7",
x"f3",
x"f4",
x"e2",
x"d4",
x"d2",
x"eb",
x"f2",
x"2c",
x"d2",
x"cb",
x"19",
x"ce",
x"dd",
x"c8",
x"ce",
x"d0",
x"d7",
x"3d",
x"b0",
x"97",
x"ee",
x"d8",
x"08",
x"18",
x"c3",
x"a1",
x"aa",
x"0b",
x"bd",
x"d1",
x"e6",
x"e2",
x"f5",
x"0b",
x"f5",
x"f4",
x"f3",
x"0f",
x"15",
x"e8",
x"00",
x"af",
x"18",
x"fc",
x"f0",
x"e2",
x"fa",
x"1d",
x"01",
x"fe",
x"fe",
x"cb",
x"25",
x"0a",
x"f1",
x"fa",
x"ec",
x"09",
x"0d",
x"05",
x"fe",
x"ef",
x"fc",
x"ff",
x"f2",
x"1a",
x"f4",
x"08",
x"19",
x"06",
x"fb",
x"f4",
x"0b",
x"f4",
x"f5",
x"15",
x"00",
x"fc",
x"0c",
x"0a",
x"02",
x"eb",
x"fe",
x"da",
x"03",
x"1b",
x"f9",
x"06",
x"11",
x"01",
x"ff",
x"f7",
x"01",
x"db",
x"00",
x"13",
x"f7",
x"fb",
x"14",
x"02",
x"fe",
x"06",
x"05",
x"d9",
x"ff",
x"1f",
x"f2",
x"01",
x"0b",
x"08",
x"fc",
x"00",
x"f7",
x"e7",
x"0d",
x"22",
x"f5",
x"f6",
x"0c",
x"fb",
x"f9",
x"11",
x"f7",
x"05",
x"e7",
x"14",
x"fa",
x"25",
x"04",
x"ed",
x"02",
x"29",
x"ff",
x"0f",
x"bc",
x"01",
x"f1",
x"1b",
x"e8",
x"fa",
x"f8",
x"37",
x"f2",
x"0e",
x"ec",
x"f1",
x"e6",
x"1b",
x"d9",
x"ec",
x"0a",
x"1b",
x"fb",
x"0f",
x"fe",
x"e9",
x"de",
x"29",
x"e3",
x"ee",
x"1d",
x"0a",
x"11",
x"12",
x"00",
x"d9",
x"df",
x"18",
x"f7",
x"f7",
x"1c",
x"ee",
x"06",
x"06",
x"05",
x"e2",
x"da",
x"16",
x"fd",
x"01",
x"f9",
x"ef",
x"f8",
x"05",
x"03",
x"df",
x"df",
x"17",
x"0e",
x"fa",
x"16",
x"dd",
x"fc",
x"13",
x"f9",
x"df",
x"f6",
x"12",
x"ff",
x"fc",
x"03",
x"02",
x"00",
x"14",
x"ff",
x"ee",
x"e6",
x"0d",
x"12",
x"ef",
x"18",
x"e8",
x"f7",
x"23",
x"0c",
x"05",
x"e6",
x"1a",
x"10",
x"fc",
x"19",
x"c8",
x"fd",
x"0a",
x"dd",
x"26",
x"fc",
x"00",
x"16",
x"eb",
x"f9",
x"85",
x"cb",
x"54",
x"e3",
x"79",
x"f4",
x"f3",
x"f2",
x"c9",
x"9a",
x"ea",
x"e3",
x"f3",
x"e1",
x"b9",
x"ad",
x"0a",
x"d0",
x"e4",
x"a1",
x"d9",
x"f1",
x"c4",
x"b4",
x"79",
x"a9",
x"00",
x"d6",
x"ad",
x"ec",
x"07",
x"e4",
x"e4",
x"d1",
x"fb",
x"e4",
x"26",
x"fa",
x"e0",
x"f0",
x"ed",
x"f5",
x"d9",
x"ea",
x"fb",
x"fd",
x"28",
x"e8",
x"e1",
x"21",
x"ff",
x"d0",
x"de",
x"d0",
x"db",
x"ee",
x"3a",
x"cc",
x"ba",
x"c7",
x"ec",
x"b1",
x"c7",
x"c5",
x"c9",
x"e1",
x"44",
x"98",
x"b6",
x"00",
x"ce",
x"cc",
x"26",
x"f4",
x"a5",
x"b3",
x"28",
x"d4",
x"c4",
x"d9",
x"ee",
x"fc",
x"10",
x"e0",
x"00",
x"01",
x"19",
x"f4",
x"f1",
x"ee",
x"e4",
x"1d",
x"e8",
x"ef",
x"02",
x"0c",
x"03",
x"08",
x"0e",
x"00",
x"c7",
x"fa",
x"f4",
x"fe",
x"1a",
x"fe",
x"f4",
x"13",
x"07",
x"0b",
x"d6",
x"e1",
x"d8",
x"00",
x"05",
x"05",
x"03",
x"18",
x"0b",
x"00",
x"ee",
x"de",
x"d4",
x"09",
x"0e",
x"fa",
x"ed",
x"18",
x"1e",
x"ed",
x"e0",
x"dc",
x"e7",
x"10",
x"10",
x"00",
x"04",
x"13",
x"0d",
x"f8",
x"f4",
x"c6",
x"dc",
x"0c",
x"09",
x"fd",
x"08",
x"0c",
x"0c",
x"03",
x"f7",
x"ca",
x"ef",
x"07",
x"0f",
x"f7",
x"0a",
x"0d",
x"16",
x"f7",
x"f8",
x"d0",
x"01",
x"19",
x"14",
x"0b",
x"00",
x"13",
x"fe",
x"00",
x"1f",
x"c8",
x"0a",
x"d0",
x"1a",
x"0f",
x"13",
x"1a",
x"fb",
x"e0",
x"32",
x"ca",
x"0a",
x"bc",
x"04",
x"ec",
x"0b",
x"07",
x"ec",
x"e5",
x"3d",
x"eb",
x"15",
x"11",
x"f9",
x"db",
x"27",
x"fb",
x"07",
x"e5",
x"0f",
x"fd",
x"0b",
x"17",
x"fb",
x"fe",
x"1b",
x"f3",
x"04",
x"08",
x"ff",
x"f3",
x"0a",
x"04",
x"f3",
x"e6",
x"19",
x"fc",
x"10",
x"fd",
x"0b",
x"fb",
x"0f",
x"f7",
x"f3",
x"f2",
x"16",
x"ff",
x"04",
x"0a",
x"f1",
x"0a",
x"0e",
x"06",
x"e0",
x"f2",
x"04",
x"01",
x"0a",
x"06",
x"f3",
x"f5",
x"0e",
x"ea",
x"bf",
x"ee",
x"0e",
x"fc",
x"1d",
x"13",
x"f9",
x"fd",
x"e8",
x"ed",
x"ae",
x"f5",
x"0b",
x"04",
x"16",
x"0c",
x"f0",
x"fc",
x"ea",
x"f1",
x"a5",
x"fc",
x"0b",
x"13",
x"10",
x"10",
x"ed",
x"eb",
x"e6",
x"cf",
x"e4",
x"13",
x"f0",
x"16",
x"f3",
x"0a",
x"a6",
x"e8",
x"78",
x"ba",
x"2a",
x"ff",
x"c9",
x"28",
x"d4",
x"be",
x"f7",
x"18",
x"0e",
x"c6",
x"a2",
x"c3",
x"ce",
x"e8",
x"c6",
x"a7",
x"e4",
x"ff",
x"ca",
x"cc",
x"6b",
x"ad",
x"ca",
x"18",
x"be",
x"f2",
x"16",
x"d6",
x"ed",
x"d4",
x"08",
x"e9",
x"0e",
x"f7",
x"da",
x"f5",
x"f7",
x"ec",
x"f5",
x"05",
x"ee",
x"08",
x"13",
x"e5",
x"df",
x"f4",
x"e2",
x"ea",
x"cb",
x"e4",
x"e2",
x"d0",
x"31",
x"d7",
x"bc",
x"c4",
x"d6",
x"d4",
x"b2",
x"d1",
x"ce",
x"c8",
x"5a",
x"ac",
x"b1",
x"03",
x"f7",
x"c8",
x"ff",
x"de",
x"de",
x"c9",
x"2e",
x"00",
x"d8",
x"de",
x"07",
x"f1",
x"ec",
x"df",
x"f5",
x"f5",
x"29",
x"f3",
x"07",
x"06",
x"f0",
x"e1",
x"e6",
x"f6",
x"04",
x"f1",
x"13",
x"1c",
x"17",
x"0a",
x"08",
x"af",
x"db",
x"ff",
x"1e",
x"0a",
x"f8",
x"14",
x"1a",
x"fe",
x"0a",
x"ae",
x"e4",
x"0e",
x"13",
x"ff",
x"17",
x"0d",
x"0a",
x"fb",
x"ec",
x"c5",
x"e3",
x"0d",
x"07",
x"09",
x"13",
x"fb",
x"0b",
x"ff",
x"05",
x"c9",
x"f9",
x"12",
x"fe",
x"0f",
x"fb",
x"0a",
x"11",
x"ff",
x"e1",
x"d2",
x"fe",
x"1e",
x"09",
x"00",
x"ec",
x"f6",
x"10",
x"00",
x"e1",
x"cc",
x"fd",
x"2a",
x"1a",
x"09",
x"fb",
x"fb",
x"06",
x"08",
x"f5",
x"d1",
x"12",
x"3d",
x"1a",
x"16",
x"dc",
x"12",
x"fd",
x"fe",
x"16",
x"d7",
x"0b",
x"f7",
x"1d",
x"06",
x"c2",
x"12",
x"00",
x"cf",
x"3b",
x"c7",
x"0d",
x"d4",
x"fb",
x"ec",
x"e8",
x"02",
x"12",
x"c8",
x"2e",
x"e2",
x"12",
x"12",
x"fd",
x"f0",
x"10",
x"04",
x"13",
x"dd",
x"10",
x"ee",
x"0f",
x"1c",
x"ee",
x"fb",
x"1f",
x"07",
x"11",
x"01",
x"00",
x"eb",
x"06",
x"01",
x"e2",
x"fd",
x"15",
x"fe",
x"0c",
x"00",
x"ff",
x"f4",
x"03",
x"00",
x"ef",
x"02",
x"11",
x"02",
x"15",
x"07",
x"e3",
x"04",
x"fb",
x"fe",
x"e4",
x"ea",
x"fb",
x"15",
x"1b",
x"0d",
x"f3",
x"03",
x"fa",
x"ff",
x"e4",
x"ee",
x"f5",
x"1a",
x"10",
x"0b",
x"09",
x"03",
x"cb",
x"09",
x"b8",
x"14",
x"fe",
x"1b",
x"17",
x"15",
x"03",
x"ed",
x"bc",
x"01",
x"75",
x"12",
x"06",
x"16",
x"1e",
x"11",
x"04",
x"bf",
x"9e",
x"e8",
x"3d",
x"25",
x"dd",
x"20",
x"22",
x"15",
x"c8",
x"00",
x"86",
x"f7",
x"46",
x"0b",
x"c7",
x"36",
x"c8",
x"df",
x"d2",
x"36",
x"1a",
x"e2",
x"01",
x"e4",
x"08",
x"06",
x"79",
x"b2",
x"cb",
x"3a",
x"dc",
x"d0",
x"4d",
x"a0",
x"0b",
x"f7",
x"bc",
x"f9",
x"07",
x"04",
x"e2",
x"d1",
x"c7",
x"e4",
x"0d",
x"d7",
x"e0",
x"00",
x"07",
x"f7",
x"f5",
x"f8",
x"f6",
x"ed",
x"ee",
x"ee",
x"ec",
x"0f",
x"df",
x"e5",
x"df",
x"0b",
x"d3",
x"e5",
x"29",
x"d6",
x"bb",
x"e7",
x"cf",
x"e6",
x"b6",
x"d3",
x"c2",
x"eb",
x"4a",
x"b9",
x"ca",
x"fb",
x"1d",
x"d5",
x"ef",
x"cb",
x"0a",
x"c3",
x"26",
x"09",
x"f1",
x"ff",
x"00",
x"b5",
x"e4",
x"ea",
x"11",
x"f1",
x"1d",
x"f6",
x"1b",
x"fb",
x"f1",
x"ae",
x"ed",
x"09",
x"23",
x"07",
x"05",
x"08",
x"15",
x"1e",
x"04",
x"ac",
x"f7",
x"15",
x"04",
x"23",
x"f9",
x"00",
x"11",
x"14",
x"00",
x"c1",
x"ea",
x"13",
x"06",
x"0a",
x"fe",
x"01",
x"0e",
x"0f",
x"0f",
x"e0",
x"f3",
x"1a",
x"fe",
x"02",
x"f0",
x"fb",
x"0e",
x"07",
x"ef",
x"f3",
x"f8",
x"17",
x"09",
x"08",
x"ea",
x"fe",
x"04",
x"07",
x"c2",
x"f7",
x"f2",
x"28",
x"0d",
x"14",
x"00",
x"e4",
x"08",
x"fe",
x"d7",
x"f8",
x"f5",
x"30",
x"19",
x"10",
x"ef",
x"00",
x"03",
x"00",
x"f6",
x"01",
x"14",
x"27",
x"1d",
x"10",
x"bf",
x"23",
x"00",
x"d8",
x"1d",
x"fd",
x"0c",
x"e7",
x"09",
x"00",
x"a6",
x"11",
x"05",
x"d5",
x"36",
x"ef",
x"05",
x"f6",
x"f6",
x"e8",
x"e3",
x"f2",
x"0a",
x"c7",
x"21",
x"e6",
x"fd",
x"0f",
x"ee",
x"08",
x"00",
x"0d",
x"17",
x"d3",
x"13",
x"f2",
x"12",
x"10",
x"e0",
x"00",
x"06",
x"15",
x"12",
x"01",
x"10",
x"fb",
x"06",
x"1a",
x"e6",
x"f9",
x"08",
x"f6",
x"12",
x"fd",
x"f4",
x"f2",
x"03",
x"04",
x"f0",
x"f3",
x"f7",
x"00",
x"09",
x"f3",
x"dc",
x"f5",
x"f0",
x"02",
x"00",
x"01",
x"f5",
x"02",
x"19",
x"fa",
x"f3",
x"f0",
x"e5",
x"10",
x"07",
x"02",
x"0c",
x"08",
x"11",
x"07",
x"f9",
x"f7",
x"d3",
x"19",
x"f8",
x"0a",
x"00",
x"fe",
x"12",
x"0c",
x"c7",
x"e6",
x"af",
x"f8",
x"d5",
x"10",
x"00",
x"00",
x"10",
x"10",
x"cc",
x"e5",
x"d2",
x"e3",
x"7f",
x"36",
x"ee",
x"fc",
x"e3",
x"04",
x"ae",
x"12",
x"db",
x"da",
x"54",
x"09",
x"fc",
x"f3",
x"b0",
x"fa",
x"ce",
x"4b",
x"fe",
x"fb",
x"ac",
x"de",
x"11",
x"02",
x"98",
x"cd",
x"cf",
x"6e",
x"cc",
x"e2",
x"26",
x"9d",
x"ed",
x"eb",
x"d3",
x"d6",
x"f2",
x"25",
x"ec",
x"db",
x"e7",
x"d7",
x"d5",
x"dc",
x"ee",
x"fb",
x"01",
x"ed",
x"e1",
x"e0",
x"1d",
x"e2",
x"f3",
x"de",
x"e1",
x"ee",
x"e8",
x"ea",
x"16",
x"0d",
x"e3",
x"ef",
x"1e",
x"ea",
x"f1",
x"d4",
x"15",
x"de",
x"e5",
x"eb",
x"be",
x"ea",
x"3d",
x"c8",
x"ca",
x"c2",
x"28",
x"e6",
x"0f",
x"00",
x"00",
x"d2",
x"00",
x"cf",
x"ff",
x"f4",
x"23",
x"cb",
x"e3",
x"1a",
x"12",
x"ca",
x"f5",
x"d3",
x"ff",
x"1f",
x"fd",
x"c4",
x"e9",
x"0f",
x"fe",
x"fa",
x"08",
x"ef",
x"08",
x"0d",
x"d6",
x"e2",
x"da",
x"17",
x"f2",
x"0a",
x"ef",
x"e3",
x"02",
x"1d",
x"ca",
x"00",
x"e8",
x"16",
x"fa",
x"0c",
x"f8",
x"d2",
x"05",
x"18",
x"00",
x"fc",
x"ff",
x"18",
x"03",
x"15",
x"f2",
x"db",
x"00",
x"0a",
x"ee",
x"fa",
x"f9",
x"0c",
x"0a",
x"13",
x"f3",
x"dc",
x"06",
x"0c",
x"c8",
x"f7",
x"f0",
x"15",
x"15",
x"0f",
x"ef",
x"f3",
x"06",
x"07",
x"d9",
x"08",
x"f9",
x"25",
x"07",
x"1c",
x"e4",
x"1d",
x"06",
x"0f",
x"fc",
x"0d",
x"1d",
x"19",
x"0e",
x"12",
x"cb",
x"1c",
x"0f",
x"f3",
x"17",
x"f8",
x"00",
x"e5",
x"01",
x"f6",
x"c9",
x"04",
x"fe",
x"b9",
x"2d",
x"02",
x"f9",
x"f7",
x"f2",
x"00",
x"e6",
x"01",
x"fc",
x"bd",
x"1b",
x"ef",
x"ff",
x"09",
x"f9",
x"ff",
x"f0",
x"fd",
x"09",
x"d2",
x"0a",
x"03",
x"09",
x"18",
x"f6",
x"0b",
x"00",
x"10",
x"14",
x"fd",
x"07",
x"f9",
x"fb",
x"24",
x"e8",
x"f1",
x"00",
x"fa",
x"0b",
x"f7",
x"d5",
x"f4",
x"f4",
x"0c",
x"fd",
x"f4",
x"17",
x"ed",
x"fe",
x"f4",
x"e0",
x"f7",
x"f5",
x"14",
x"ec",
x"fe",
x"1d",
x"f3",
x"f7",
x"04",
x"f1",
x"fe",
x"ec",
x"11",
x"01",
x"03",
x"15",
x"ee",
x"04",
x"08",
x"e7",
x"ec",
x"fd",
x"00",
x"f9",
x"ff",
x"0f",
x"fa",
x"08",
x"10",
x"03",
x"f1",
x"f6",
x"fc",
x"11",
x"1a",
x"19",
x"dc",
x"f6",
x"08",
x"f3",
x"f4",
x"00",
x"f2",
x"ef",
x"0d",
x"20",
x"c5",
x"cd",
x"11",
x"00",
x"06",
x"f5",
x"d6",
x"d8",
x"f9",
x"f4",
x"d4",
x"8e",
x"06",
x"f8",
x"2f",
x"b8",
x"e0",
x"a4",
x"ff",
x"f3",
x"09",
x"c2",
x"c0",
x"01",
x"6c",
x"d2",
x"b3",
x"b9",
x"b0",
x"c9",
x"db",
x"e5",
x"e2",
x"f4",
x"3a",
x"dc",
x"dd",
x"de",
x"d8",
x"dc",
x"e2",
x"e8",
x"ea",
x"fa",
x"fe",
x"ea",
x"f2",
x"11",
x"e6",
x"1c",
x"e0",
x"ea",
x"f6",
x"06",
x"e8",
x"1d",
x"23",
x"fc",
x"07",
x"f5",
x"fb",
x"f8",
x"e0",
x"22",
x"e4",
x"14",
x"1c",
x"bd",
x"ee",
x"13",
x"db",
x"af",
x"bd",
x"26",
x"0d",
x"fa",
x"fc",
x"ef",
x"bb",
x"11",
x"e3",
x"eb",
x"11",
x"0a",
x"0a",
x"f7",
x"1b",
x"05",
x"b0",
x"f0",
x"b9",
x"0b",
x"13",
x"d3",
x"1e",
x"f8",
x"04",
x"e2",
x"e1",
x"f1",
x"c4",
x"01",
x"04",
x"cc",
x"14",
x"fd",
x"0c",
x"dc",
x"02",
x"f3",
x"c4",
x"ee",
x"1e",
x"f7",
x"00",
x"ec",
x"15",
x"e6",
x"0f",
x"e9",
x"d9",
x"00",
x"16",
x"ff",
x"fd",
x"e4",
x"15",
x"01",
x"fe",
x"e0",
x"e5",
x"03",
x"18",
x"ee",
x"01",
x"fb",
x"18",
x"0b",
x"0c",
x"ed",
x"fb",
x"fd",
x"12",
x"d3",
x"06",
x"f4",
x"13",
x"0e",
x"12",
x"f0",
x"03",
x"01",
x"00",
x"fe",
x"07",
x"03",
x"15",
x"09",
x"1d",
x"e2",
x"05",
x"12",
x"04",
x"09",
x"02",
x"0f",
x"18",
x"0e",
x"0b",
x"e1",
x"13",
x"08",
x"c5",
x"24",
x"05",
x"fa",
x"f1",
x"f1",
x"f3",
x"d6",
x"0a",
x"fa",
x"bc",
x"27",
x"f5",
x"f9",
x"07",
x"e8",
x"14",
x"eb",
x"03",
x"ee",
x"d8",
x"0c",
x"01",
x"0b",
x"18",
x"e6",
x"02",
x"03",
x"00",
x"00",
x"e4",
x"0c",
x"05",
x"00",
x"1f",
x"f6",
x"00",
x"f9",
x"04",
x"10",
x"e9",
x"e7",
x"f5",
x"ec",
x"17",
x"ef",
x"f9",
x"1e",
x"ec",
x"05",
x"f1",
x"cb",
x"f5",
x"fc",
x"00",
x"04",
x"f6",
x"19",
x"ed",
x"fe",
x"fb",
x"bd",
x"06",
x"00",
x"12",
x"f2",
x"fd",
x"0e",
x"ef",
x"fe",
x"0b",
x"de",
x"ec",
x"11",
x"f4",
x"fd",
x"07",
x"20",
x"e7",
x"01",
x"02",
x"e1",
x"f8",
x"10",
x"fa",
x"f7",
x"12",
x"1a",
x"dd",
x"f0",
x"03",
x"e5",
x"e5",
x"1e",
x"0f",
x"f8",
x"03",
x"23",
x"eb",
x"fa",
x"12",
x"cb",
x"e3",
x"22",
x"ff",
x"0b",
x"fb",
x"12",
x"df",
x"eb",
x"11",
x"e3",
x"01",
x"02",
x"c0",
x"0b",
x"f8",
x"e8",
x"cb",
x"98",
x"f7",
x"e7",
x"30",
x"8c",
x"d2",
x"d1",
x"0c",
x"b5",
x"f2",
x"c6",
x"b4",
x"f0",
x"5f",
x"01",
x"06",
x"b1",
x"a9",
x"d6",
x"ac",
x"ea",
x"d4",
x"da",
x"33",
x"e9",
x"e2",
x"de",
x"df",
x"e8",
x"e2",
x"cd",
x"ee",
x"04",
x"04",
x"f3",
x"f3",
x"eb",
x"f8",
x"14",
x"ec",
x"f5",
x"f4",
x"0b",
x"ee",
x"1b",
x"00",
x"f4",
x"f8",
x"ec",
x"e7",
x"f2",
x"e9",
x"29",
x"e6",
x"37",
x"f6",
x"a1",
x"f5",
x"e7",
x"e1",
x"c4",
x"d0",
x"e9",
x"18",
x"0d",
x"ee",
x"01",
x"c5",
x"f9",
x"12",
x"f1",
x"03",
x"f0",
x"1a",
x"0d",
x"db",
x"fd",
x"d5",
x"f7",
x"d2",
x"0c",
x"13",
x"e8",
x"16",
x"07",
x"ff",
x"f2",
x"f6",
x"f1",
x"e5",
x"ff",
x"00",
x"f1",
x"1f",
x"ef",
x"03",
x"ef",
x"0a",
x"05",
x"ee",
x"f2",
x"0f",
x"f3",
x"ff",
x"ee",
x"1f",
x"d7",
x"0e",
x"09",
x"f9",
x"fb",
x"11",
x"ec",
x"f8",
x"de",
x"1a",
x"df",
x"0c",
x"00",
x"fd",
x"0d",
x"11",
x"00",
x"fd",
x"f2",
x"16",
x"f8",
x"16",
x"ef",
x"00",
x"02",
x"12",
x"f5",
x"08",
x"f5",
x"05",
x"f0",
x"0a",
x"e4",
x"02",
x"10",
x"04",
x"eb",
x"0e",
x"02",
x"03",
x"00",
x"2c",
x"d6",
x"09",
x"0f",
x"eb",
x"f3",
x"11",
x"0c",
x"00",
x"0a",
x"f2",
x"f1",
x"13",
x"06",
x"ae",
x"12",
x"15",
x"08",
x"06",
x"f7",
x"fa",
x"f5",
x"04",
x"ec",
x"be",
x"31",
x"f8",
x"f0",
x"0f",
x"ef",
x"04",
x"e6",
x"ee",
x"eb",
x"e0",
x"ff",
x"00",
x"ec",
x"26",
x"f9",
x"00",
x"06",
x"05",
x"ff",
x"e7",
x"00",
x"15",
x"f0",
x"1d",
x"ef",
x"f4",
x"fa",
x"03",
x"0a",
x"fc",
x"cb",
x"07",
x"f6",
x"07",
x"ec",
x"f0",
x"13",
x"ee",
x"fb",
x"fc",
x"d1",
x"f8",
x"0c",
x"12",
x"ff",
x"ff",
x"09",
x"ea",
x"00",
x"fd",
x"d0",
x"00",
x"11",
x"06",
x"01",
x"03",
x"10",
x"ea",
x"ec",
x"0f",
x"ee",
x"fe",
x"10",
x"14",
x"f8",
x"09",
x"10",
x"ee",
x"fc",
x"08",
x"f8",
x"10",
x"14",
x"15",
x"f4",
x"00",
x"0b",
x"e9",
x"da",
x"00",
x"f0",
x"0a",
x"12",
x"fe",
x"05",
x"fc",
x"02",
x"ea",
x"07",
x"06",
x"cd",
x"08",
x"19",
x"f7",
x"0e",
x"f3",
x"f0",
x"06",
x"e4",
x"f3",
x"f8",
x"13",
x"2d",
x"d6",
x"13",
x"00",
x"e8",
x"f4",
x"9a",
x"ca",
x"b8",
x"4c",
x"4b",
x"c4",
x"d1",
x"f0",
x"8e",
x"c3",
x"9b",
x"b6",
x"e7",
x"70",
x"ad",
x"da",
x"94",
x"94",
x"b0",
x"97",
x"de",
x"fc",
x"dc",
x"29",
x"d0",
x"d0",
x"db",
x"d5",
x"dd",
x"e4",
x"c4",
x"fd",
x"fa",
x"f6",
x"fa",
x"03",
x"f9",
x"fd",
x"fc",
x"f7",
x"fa",
x"f8",
x"23",
x"e0",
x"28",
x"f7",
x"e7",
x"e9",
x"e6",
x"dd",
x"e1",
x"c7",
x"05",
x"f1",
x"23",
x"14",
x"b4",
x"e7",
x"f2",
x"d9",
x"c8",
x"c2",
x"f2",
x"12",
x"26",
x"c7",
x"fa",
x"cc",
x"f7",
x"e4",
x"f3",
x"08",
x"08",
x"14",
x"10",
x"df",
x"00",
x"c2",
x"0c",
x"ec",
x"ea",
x"0f",
x"dc",
x"14",
x"03",
x"f7",
x"0c",
x"fb",
x"06",
x"e0",
x"f8",
x"15",
x"d6",
x"16",
x"00",
x"00",
x"1e",
x"fd",
x"02",
x"f5",
x"fa",
x"0d",
x"f6",
x"07",
x"01",
x"0f",
x"f4",
x"07",
x"f0",
x"10",
x"09",
x"0c",
x"fd",
x"0b",
x"f5",
x"14",
x"dd",
x"16",
x"f1",
x"12",
x"fe",
x"10",
x"f2",
x"0f",
x"da",
x"08",
x"d8",
x"0b",
x"ec",
x"17",
x"05",
x"1d",
x"fa",
x"0c",
x"c8",
x"fa",
x"db",
x"1e",
x"d9",
x"04",
x"05",
x"00",
x"e1",
x"0a",
x"d3",
x"f0",
x"db",
x"25",
x"e9",
x"0e",
x"04",
x"f8",
x"03",
x"17",
x"e4",
x"02",
x"d8",
x"0c",
x"fb",
x"22",
x"0a",
x"c1",
x"19",
x"12",
x"e5",
x"12",
x"dd",
x"00",
x"06",
x"00",
x"f1",
x"d3",
x"28",
x"07",
x"dc",
x"21",
x"de",
x"0f",
x"fc",
x"00",
x"f5",
x"e6",
x"00",
x"19",
x"eb",
x"16",
x"f1",
x"f3",
x"01",
x"f9",
x"00",
x"f6",
x"ea",
x"00",
x"f7",
x"11",
x"fb",
x"fb",
x"f9",
x"00",
x"ff",
x"01",
x"ca",
x"02",
x"10",
x"15",
x"0c",
x"fb",
x"fc",
x"f5",
x"00",
x"ff",
x"e8",
x"04",
x"0a",
x"0f",
x"09",
x"09",
x"11",
x"f0",
x"00",
x"fd",
x"ff",
x"f8",
x"1d",
x"03",
x"fe",
x"06",
x"03",
x"f5",
x"f8",
x"05",
x"fa",
x"fc",
x"09",
x"fd",
x"03",
x"09",
x"0b",
x"f9",
x"fc",
x"fb",
x"02",
x"ff",
x"08",
x"0f",
x"06",
x"f9",
x"fe",
x"f7",
x"fd",
x"0e",
x"00",
x"01",
x"13",
x"fa",
x"fd",
x"06",
x"07",
x"f5",
x"f1",
x"f5",
x"eb",
x"05",
x"18",
x"02",
x"0d",
x"09",
x"f8",
x"0c",
x"e2",
x"fd",
x"04",
x"12",
x"f5",
x"da",
x"19",
x"f7",
x"05",
x"17",
x"91",
x"e5",
x"da",
x"52",
x"6a",
x"ab",
x"b9",
x"e6",
x"01",
x"87",
x"da",
x"be",
x"e6",
x"50",
x"b9",
x"d2",
x"a2",
x"99",
x"0b",
x"a7",
x"cd",
x"1f",
x"d2",
x"41",
x"d9",
x"cc",
x"c7",
x"c5",
x"cf",
x"d7",
x"d4",
x"e2",
x"f2",
x"e5",
x"d5",
x"e9",
x"db",
x"f4",
x"22",
x"dd",
x"14",
x"fc",
x"17",
x"dd",
x"26",
x"00",
x"ea",
x"fd",
x"04",
x"d6",
x"e9",
x"bf",
x"e5",
x"e1",
x"0f",
x"03",
x"c2",
x"e4",
x"22",
x"c0",
x"cc",
x"a2",
x"d2",
x"f3",
x"42",
x"f0",
x"f1",
x"da",
x"f2",
x"8c",
x"d6",
x"f6",
x"ab",
x"12",
x"0c",
x"df",
x"19",
x"dc",
x"0b",
x"e4",
x"df",
x"f6",
x"bc",
x"19",
x"01",
x"f2",
x"18",
x"e8",
x"04",
x"e6",
x"e4",
x"fe",
x"b2",
x"16",
x"00",
x"ff",
x"29",
x"f3",
x"d6",
x"f1",
x"01",
x"0f",
x"e4",
x"1f",
x"fc",
x"0f",
x"10",
x"0c",
x"e3",
x"02",
x"07",
x"12",
x"02",
x"0b",
x"f9",
x"06",
x"f4",
x"0c",
x"f0",
x"12",
x"fb",
x"13",
x"f9",
x"02",
x"e0",
x"0d",
x"eb",
x"12",
x"e9",
x"11",
x"09",
x"13",
x"e8",
x"0a",
x"d1",
x"e4",
x"d9",
x"1d",
x"df",
x"18",
x"12",
x"07",
x"e9",
x"02",
x"d6",
x"f8",
x"e1",
x"0f",
x"fa",
x"15",
x"0b",
x"ee",
x"01",
x"17",
x"d0",
x"0c",
x"f3",
x"24",
x"04",
x"13",
x"f5",
x"ca",
x"0c",
x"0c",
x"cc",
x"2c",
x"06",
x"18",
x"05",
x"fd",
x"f6",
x"e1",
x"14",
x"11",
x"de",
x"18",
x"08",
x"00",
x"01",
x"ef",
x"00",
x"ed",
x"f3",
x"03",
x"09",
x"0c",
x"00",
x"08",
x"f9",
x"f8",
x"07",
x"ee",
x"dc",
x"13",
x"1b",
x"0c",
x"08",
x"12",
x"f2",
x"f1",
x"f4",
x"f5",
x"e6",
x"0b",
x"15",
x"ea",
x"0d",
x"09",
x"00",
x"f8",
x"00",
x"f5",
x"fa",
x"05",
x"02",
x"f1",
x"f6",
x"12",
x"ff",
x"fa",
x"f9",
x"f4",
x"fc",
x"03",
x"11",
x"00",
x"fc",
x"00",
x"f7",
x"00",
x"ff",
x"f8",
x"0d",
x"01",
x"00",
x"00",
x"0e",
x"00",
x"f3",
x"f9",
x"02",
x"f6",
x"0a",
x"02",
x"0e",
x"fb",
x"04",
x"04",
x"f6",
x"fb",
x"f0",
x"07",
x"e8",
x"11",
x"21",
x"e1",
x"07",
x"f7",
x"f0",
x"0d",
x"ed",
x"fd",
x"ea",
x"15",
x"06",
x"e4",
x"0e",
x"01",
x"cc",
x"f0",
x"df",
x"e3",
x"f8",
x"38",
x"ca",
x"da",
x"06",
x"de",
x"dd",
x"e0",
x"a5",
x"d5",
x"f5",
x"44",
x"58",
x"a7",
x"c7",
x"f9",
x"f5",
x"8c",
x"e6",
x"cc",
x"ff",
x"1c",
x"c0",
x"db",
x"c8",
x"d3",
x"18",
x"af",
x"b4",
x"df",
x"27",
x"26",
x"de",
x"fb",
x"e5",
x"d9",
x"e6",
x"dc",
x"cb",
x"03",
x"16",
x"f9",
x"f6",
x"06",
x"ff",
x"f3",
x"f6",
x"e7",
x"f9",
x"1e",
x"fd",
x"ca",
x"e4",
x"cc",
x"e7",
x"df",
x"19",
x"d7",
x"be",
x"fc",
x"f1",
x"d8",
x"f7",
x"fe",
x"0b",
x"d9",
x"19",
x"b7",
x"be",
x"cb",
x"d4",
x"d8",
x"38",
x"1a",
x"e7",
x"cc",
x"03",
x"c2",
x"d6",
x"f6",
x"a1",
x"06",
x"0a",
x"fb",
x"12",
x"f7",
x"fe",
x"e0",
x"c5",
x"fd",
x"8c",
x"01",
x"1e",
x"0a",
x"ff",
x"f1",
x"e1",
x"04",
x"e8",
x"00",
x"db",
x"06",
x"01",
x"00",
x"15",
x"f5",
x"ce",
x"f6",
x"ef",
x"04",
x"f7",
x"13",
x"f8",
x"eb",
x"0c",
x"fe",
x"d4",
x"f6",
x"08",
x"10",
x"f8",
x"11",
x"fe",
x"ef",
x"1b",
x"04",
x"e6",
x"07",
x"f6",
x"ff",
x"05",
x"12",
x"ff",
x"e2",
x"08",
x"0b",
x"ee",
x"0e",
x"e5",
x"18",
x"f5",
x"15",
x"f4",
x"df",
x"00",
x"23",
x"ea",
x"09",
x"fd",
x"11",
x"ee",
x"12",
x"ec",
x"f2",
x"09",
x"2a",
x"fd",
x"04",
x"fd",
x"0b",
x"f8",
x"0a",
x"f2",
x"e5",
x"0b",
x"22",
x"02",
x"fc",
x"00",
x"ed",
x"06",
x"13",
x"e9",
x"f6",
x"04",
x"00",
x"07",
x"ea",
x"f4",
x"ed",
x"f4",
x"0f",
x"ec",
x"0c",
x"00",
x"08",
x"09",
x"ea",
x"f1",
x"f3",
x"fc",
x"06",
x"fc",
x"06",
x"0c",
x"16",
x"f4",
x"fa",
x"f0",
x"f6",
x"00",
x"0b",
x"0a",
x"fa",
x"f8",
x"10",
x"e6",
x"00",
x"01",
x"fc",
x"f7",
x"02",
x"0a",
x"f8",
x"fe",
x"09",
x"ee",
x"fd",
x"f5",
x"fe",
x"05",
x"00",
x"15",
x"f9",
x"09",
x"0c",
x"d9",
x"fe",
x"ee",
x"ee",
x"10",
x"fe",
x"05",
x"f2",
x"00",
x"f9",
x"e8",
x"fc",
x"fd",
x"fc",
x"08",
x"02",
x"03",
x"ec",
x"ff",
x"00",
x"ef",
x"00",
x"fe",
x"00",
x"fd",
x"07",
x"13",
x"fb",
x"fb",
x"00",
x"e7",
x"f8",
x"f4",
x"11",
x"e5",
x"06",
x"f7",
x"cf",
x"0c",
x"f9",
x"e1",
x"0b",
x"eb",
x"e7",
x"f3",
x"08",
x"fd",
x"ce",
x"fe",
x"fe",
x"bf",
x"17",
x"e8",
x"fe",
x"03",
x"1e",
x"d0",
x"cd",
x"09",
x"e2",
x"f4",
x"d7",
x"d5",
x"a8",
x"0d",
x"35",
x"6e",
x"c2",
x"de",
x"c5",
x"e7",
x"73",
x"e7",
x"d4",
x"01",
x"36",
x"d0",
x"ea",
x"bf",
x"bc",
x"d9",
x"b6",
x"d2",
x"e3",
x"1c",
x"02",
x"e3",
x"00",
x"df",
x"d6",
x"ef",
x"d5",
x"e4",
x"f9",
x"09",
x"00",
x"00",
x"07",
x"fb",
x"f6",
x"03",
x"00",
x"07",
x"11",
x"ef",
x"cc",
x"09",
x"e8",
x"e3",
x"dc",
x"16",
x"e5",
x"e2",
x"e2",
x"df",
x"02",
x"f1",
x"0c",
x"07",
x"e2",
x"f7",
x"c2",
x"d6",
x"dc",
x"e5",
x"fd",
x"33",
x"06",
x"ee",
x"bf",
x"bc",
x"b7",
x"cc",
x"02",
x"ee",
x"16",
x"0b",
x"fe",
x"fd",
x"f7",
x"bf",
x"e1",
x"f1",
x"07",
x"bf",
x"0c",
x"0c",
x"e1",
x"0b",
x"e9",
x"d5",
x"f2",
x"02",
x"fd",
x"f7",
x"09",
x"0c",
x"f3",
x"f7",
x"f1",
x"bb",
x"fc",
x"f7",
x"fb",
x"fa",
x"18",
x"06",
x"dc",
x"f4",
x"00",
x"c1",
x"05",
x"db",
x"09",
x"08",
x"10",
x"0c",
x"d5",
x"0d",
x"fb",
x"eb",
x"01",
x"e4",
x"03",
x"fc",
x"0f",
x"0a",
x"e3",
x"07",
x"0f",
x"e7",
x"f4",
x"de",
x"10",
x"09",
x"10",
x"02",
x"e1",
x"09",
x"1b",
x"e4",
x"fb",
x"cb",
x"2b",
x"12",
x"11",
x"f8",
x"f3",
x"11",
x"11",
x"ff",
x"ef",
x"e2",
x"0d",
x"06",
x"05",
x"f7",
x"ea",
x"00",
x"1e",
x"06",
x"03",
x"dd",
x"05",
x"f9",
x"f8",
x"f5",
x"e7",
x"02",
x"13",
x"fd",
x"f6",
x"f6",
x"f0",
x"03",
x"fe",
x"00",
x"fa",
x"f3",
x"16",
x"f5",
x"ea",
x"e8",
x"f7",
x"fa",
x"02",
x"f1",
x"fb",
x"f3",
x"15",
x"ef",
x"02",
x"e8",
x"ee",
x"0d",
x"00",
x"fe",
x"01",
x"07",
x"07",
x"e7",
x"fb",
x"ef",
x"ed",
x"09",
x"f7",
x"03",
x"00",
x"02",
x"04",
x"da",
x"f7",
x"eb",
x"f5",
x"24",
x"05",
x"05",
x"f7",
x"01",
x"05",
x"d1",
x"fe",
x"fa",
x"f7",
x"14",
x"0a",
x"02",
x"eb",
x"07",
x"09",
x"df",
x"fa",
x"06",
x"f6",
x"fe",
x"11",
x"08",
x"f2",
x"f9",
x"fe",
x"d0",
x"00",
x"f9",
x"fc",
x"01",
x"14",
x"01",
x"f7",
x"07",
x"00",
x"d5",
x"04",
x"df",
x"fc",
x"e7",
x"01",
x"ec",
x"e1",
x"1c",
x"e7",
x"cb",
x"0f",
x"e6",
x"eb",
x"e0",
x"11",
x"f8",
x"db",
x"12",
x"f0",
x"c0",
x"04",
x"e3",
x"e9",
x"00",
x"23",
x"cc",
x"e2",
x"f4",
x"d7",
x"f6",
x"d1",
x"05",
x"af",
x"05",
x"2c",
x"83",
x"ca",
x"ff",
x"d5",
x"fb",
x"90",
x"1c",
x"e5",
x"14",
x"0a",
x"f8",
x"dd",
x"c7",
x"f6",
x"d9",
x"b9",
x"c7",
x"f5",
x"1a",
x"e4",
x"eb",
x"e6",
x"13",
x"e9",
x"fd",
x"dc",
x"f4",
x"07",
x"25",
x"fc",
x"f1",
x"f5",
x"06",
x"fa",
x"02",
x"eb",
x"f8",
x"e8",
x"f3",
x"e7",
x"0e",
x"f3",
x"d3",
x"e5",
x"e5",
x"ea",
x"de",
x"da",
x"e4",
x"fb",
x"0e",
x"03",
x"cf",
x"e9",
x"e0",
x"cf",
x"da",
x"e8",
x"0a",
x"00",
x"12",
x"e9",
x"f2",
x"cd",
x"9f",
x"af",
x"b0",
x"f4",
x"17",
x"fb",
x"16",
x"de",
x"16",
x"d7",
x"c3",
x"dc",
x"eb",
x"00",
x"28",
x"fa",
x"02",
x"04",
x"00",
x"e1",
x"dc",
x"02",
x"fe",
x"f9",
x"13",
x"0a",
x"10",
x"cd",
x"0f",
x"de",
x"cc",
x"01",
x"e7",
x"fd",
x"07",
x"08",
x"00",
x"ca",
x"05",
x"03",
x"df",
x"10",
x"f1",
x"f5",
x"12",
x"fe",
x"06",
x"fd",
x"0b",
x"07",
x"f6",
x"f5",
x"ee",
x"03",
x"0a",
x"11",
x"f0",
x"f1",
x"0b",
x"00",
x"f2",
x"00",
x"f1",
x"12",
x"14",
x"04",
x"f7",
x"fa",
x"09",
x"0a",
x"f6",
x"f8",
x"ec",
x"18",
x"fd",
x"0e",
x"f9",
x"f7",
x"05",
x"18",
x"ef",
x"f8",
x"e5",
x"0c",
x"f9",
x"00",
x"f8",
x"e8",
x"01",
x"25",
x"fa",
x"ff",
x"ed",
x"02",
x"f4",
x"f4",
x"fe",
x"ec",
x"00",
x"25",
x"f3",
x"fd",
x"e9",
x"f6",
x"02",
x"fb",
x"f4",
x"f4",
x"00",
x"23",
x"f4",
x"02",
x"f0",
x"ff",
x"03",
x"f1",
x"04",
x"03",
x"fe",
x"1b",
x"f2",
x"f3",
x"f3",
x"fc",
x"05",
x"06",
x"08",
x"fa",
x"09",
x"0e",
x"f3",
x"fa",
x"ed",
x"e9",
x"03",
x"09",
x"fe",
x"06",
x"05",
x"19",
x"e9",
x"f6",
x"eb",
x"ec",
x"1b",
x"0b",
x"0a",
x"f8",
x"fe",
x"12",
x"e6",
x"00",
x"eb",
x"ea",
x"03",
x"1e",
x"0c",
x"01",
x"04",
x"fd",
x"e1",
x"03",
x"ed",
x"ed",
x"17",
x"07",
x"01",
x"ff",
x"13",
x"00",
x"e2",
x"07",
x"f6",
x"f9",
x"0d",
x"0d",
x"f2",
x"fe",
x"16",
x"ea",
x"df",
x"04",
x"fa",
x"02",
x"db",
x"23",
x"f4",
x"0a",
x"1c",
x"07",
x"d0",
x"16",
x"ec",
x"e4",
x"da",
x"32",
x"e5",
x"fc",
x"0d",
x"e9",
x"c1",
x"ee",
x"04",
x"da",
x"01",
x"17",
x"a4",
x"ef",
x"03",
x"e0",
x"f0",
x"af",
x"1b",
x"c0",
x"15",
x"2a",
x"a4",
x"dc",
x"0b",
x"f0",
x"1c",
x"ae",
x"12",
x"2c",
x"f8",
x"02",
x"ef",
x"d3",
x"ef",
x"1b",
x"db",
x"b1",
x"d1",
x"1b",
x"fc",
x"fc",
x"00",
x"08",
x"fa",
x"f8",
x"00",
x"f0",
x"00",
x"07",
x"23",
x"f9",
x"ea",
x"fd",
x"00",
x"07",
x"f7",
x"f8",
x"00",
x"fc",
x"fc",
x"f5",
x"0b",
x"fa",
x"e8",
x"04",
x"ee",
x"f9",
x"00",
x"c7",
x"f4",
x"f8",
x"0d",
x"e8",
x"a0",
x"00",
x"cb",
x"da",
x"c0",
x"d2",
x"fd",
x"0a",
x"05",
x"da",
x"d3",
x"dd",
x"97",
x"dd",
x"e4",
x"cb",
x"1c",
x"0b",
x"10",
x"c7",
x"03",
x"c3",
x"c7",
x"ec",
x"fc",
x"00",
x"51",
x"06",
x"fb",
x"cc",
x"00",
x"c1",
x"0d",
x"f8",
x"e0",
x"06",
x"1e",
x"1c",
x"01",
x"d8",
x"f1",
x"aa",
x"f2",
x"0e",
x"e3",
x"03",
x"00",
x"08",
x"04",
x"e7",
x"00",
x"ee",
x"0a",
x"02",
x"ed",
x"06",
x"fd",
x"12",
x"f8",
x"ef",
x"00",
x"0d",
x"02",
x"f9",
x"fc",
x"0c",
x"01",
x"0d",
x"00",
x"e3",
x"06",
x"0a",
x"ef",
x"f1",
x"00",
x"fe",
x"f0",
x"04",
x"00",
x"ee",
x"00",
x"0e",
x"ff",
x"fc",
x"05",
x"10",
x"e8",
x"07",
x"08",
x"f3",
x"0e",
x"05",
x"f4",
x"05",
x"f7",
x"06",
x"df",
x"05",
x"00",
x"f1",
x"0b",
x"07",
x"f5",
x"0e",
x"ff",
x"15",
x"e3",
x"05",
x"fd",
x"f3",
x"0c",
x"04",
x"f3",
x"0d",
x"f8",
x"03",
x"fc",
x"f3",
x"f3",
x"ec",
x"02",
x"fe",
x"f9",
x"0a",
x"fd",
x"fb",
x"02",
x"f8",
x"fb",
x"f4",
x"f9",
x"0f",
x"f9",
x"f8",
x"e5",
x"f7",
x"06",
x"00",
x"04",
x"f5",
x"08",
x"0c",
x"f7",
x"fe",
x"f6",
x"f7",
x"12",
x"02",
x"01",
x"09",
x"00",
x"07",
x"eb",
x"fe",
x"ef",
x"f6",
x"1b",
x"0f",
x"06",
x"02",
x"12",
x"01",
x"eb",
x"00",
x"f8",
x"fa",
x"12",
x"05",
x"0e",
x"0e",
x"0b",
x"06",
x"e9",
x"f6",
x"d6",
x"fe",
x"18",
x"11",
x"09",
x"ff",
x"10",
x"13",
x"dc",
x"f5",
x"f8",
x"f8",
x"00",
x"0d",
x"f5",
x"18",
x"08",
x"10",
x"d1",
x"02",
x"fb",
x"12",
x"d2",
x"1c",
x"0b",
x"01",
x"0e",
x"e5",
x"c8",
x"00",
x"04",
x"f9",
x"ed",
x"0d",
x"e8",
x"02",
x"10",
x"bf",
x"9e",
x"ef",
x"0e",
x"d4",
x"ff",
x"26",
x"8e",
x"f8",
x"10",
x"a7",
x"f9",
x"c6",
x"15",
x"ce",
x"1f",
x"11",
x"c6",
x"eb",
x"0b",
x"dc",
x"0b",
x"de",
x"00",
x"1a",
x"28",
x"e6",
x"ff",
x"24",
x"1a",
x"1a",
x"d2",
x"c7",
x"d0",
x"1b",
x"f9",
x"fc",
x"fd",
x"f7",
x"f2",
x"fb",
x"01",
x"f2",
x"03",
x"06",
x"06",
x"f9",
x"fe",
x"01",
x"00",
x"06",
x"0a",
x"02",
x"f6",
x"03",
x"04",
x"06",
x"0a",
x"fe",
x"f6",
x"06",
x"fe",
x"00",
x"fd",
x"ed",
x"d9",
x"ca",
x"31",
x"f3",
x"ed",
x"f4",
x"c4",
x"d0",
x"c0",
x"be",
x"c1",
x"e3",
x"24",
x"cf",
x"ef",
x"f0",
x"a6",
x"db",
x"f3",
x"be",
x"ce",
x"fd",
x"33",
x"a9",
x"17",
x"e8",
x"fc",
x"e1",
x"cc",
x"e7",
x"18",
x"fb",
x"1a",
x"d5",
x"28",
x"e4",
x"11",
x"db",
x"e6",
x"00",
x"22",
x"04",
x"1f",
x"05",
x"fe",
x"a6",
x"10",
x"e9",
x"e6",
x"fe",
x"00",
x"fd",
x"18",
x"fe",
x"e5",
x"c1",
x"1a",
x"eb",
x"e8",
x"f3",
x"f7",
x"f2",
x"00",
x"ff",
x"03",
x"d2",
x"e8",
x"f9",
x"06",
x"0a",
x"f4",
x"fe",
x"05",
x"fd",
x"fc",
x"e2",
x"f0",
x"f9",
x"ee",
x"0f",
x"f0",
x"e9",
x"09",
x"fb",
x"0f",
x"df",
x"f3",
x"01",
x"f4",
x"0b",
x"f5",
x"fc",
x"06",
x"f5",
x"01",
x"db",
x"e6",
x"00",
x"ee",
x"13",
x"fc",
x"fb",
x"f4",
x"ef",
x"0c",
x"eb",
x"e8",
x"0c",
x"f4",
x"0b",
x"f7",
x"f2",
x"05",
x"f3",
x"01",
x"fa",
x"e4",
x"15",
x"f0",
x"0d",
x"e9",
x"f1",
x"fc",
x"f7",
x"0b",
x"fe",
x"f0",
x"06",
x"ee",
x"01",
x"01",
x"f6",
x"f5",
x"00",
x"00",
x"f3",
x"00",
x"12",
x"e9",
x"fb",
x"0b",
x"f3",
x"e5",
x"00",
x"04",
x"f8",
x"f3",
x"09",
x"e9",
x"0b",
x"19",
x"f3",
x"ff",
x"00",
x"f4",
x"ee",
x"f4",
x"02",
x"f0",
x"e8",
x"07",
x"18",
x"11",
x"0b",
x"ed",
x"fb",
x"eb",
x"0d",
x"f1",
x"e6",
x"fd",
x"0f",
x"06",
x"0a",
x"f5",
x"fb",
x"dd",
x"f9",
x"f1",
x"dd",
x"04",
x"13",
x"03",
x"06",
x"01",
x"f5",
x"d6",
x"fe",
x"fe",
x"ed",
x"dd",
x"23",
x"ff",
x"15",
x"e9",
x"ee",
x"c4",
x"0b",
x"04",
x"00",
x"e4",
x"1a",
x"d8",
x"db",
x"f8",
x"da",
x"d3",
x"ff",
x"21",
x"e1",
x"da",
x"1b",
x"ca",
x"e6",
x"0a",
x"b0",
x"aa",
x"06",
x"25",
x"d4",
x"e6",
x"24",
x"e3",
x"dd",
x"0d",
x"cd",
x"f9",
x"e0",
x"17",
x"e9",
x"04",
x"1c",
x"e9",
x"fd",
x"0b",
x"d5",
x"fe",
x"cb",
x"f6",
x"ec",
x"19",
x"f0",
x"12",
x"27",
x"19",
x"f6",
x"e1",
x"bc",
x"e2",
x"f9",
x"f8",
x"03",
x"f9",
x"f6",
x"f9",
x"05",
x"02",
x"f9",
x"06",
x"ff",
x"06",
x"fc",
x"fa",
x"08",
x"0a",
x"ff",
x"f7",
x"fa",
x"09",
x"03",
x"f9",
x"0a",
x"f9",
x"07",
x"05",
x"fc",
x"fa",
x"02",
x"fb",
x"eb",
x"fc",
x"d9",
x"01",
x"f2",
x"da",
x"07",
x"ea",
x"e6",
x"dc",
x"dc",
x"d9",
x"ac",
x"37",
x"ee",
x"07",
x"05",
x"e2",
x"c9",
x"ae",
x"fa",
x"ba",
x"c6",
x"2b",
x"af",
x"f2",
x"fb",
x"24",
x"a9",
x"00",
x"f8",
x"03",
x"c7",
x"0c",
x"03",
x"0e",
x"f3",
x"2d",
x"c3",
x"13",
x"e0",
x"05",
x"db",
x"22",
x"15",
x"fe",
x"db",
x"27",
x"eb",
x"fd",
x"e6",
x"f5",
x"eb",
x"24",
x"fd",
x"09",
x"b9",
x"0a",
x"f4",
x"07",
x"ff",
x"e7",
x"fc",
x"07",
x"03",
x"ff",
x"9f",
x"fe",
x"08",
x"f6",
x"fb",
x"f5",
x"f3",
x"fe",
x"fc",
x"1a",
x"8d",
x"fc",
x"05",
x"ed",
x"01",
x"ed",
x"ed",
x"13",
x"f7",
x"02",
x"75",
x"f8",
x"f9",
x"f5",
x"ec",
x"d8",
x"f7",
x"05",
x"08",
x"02",
x"ab",
x"f6",
x"00",
x"e6",
x"fa",
x"e4",
x"fc",
x"fa",
x"f6",
x"00",
x"c5",
x"f4",
x"fa",
x"ec",
x"fb",
x"d8",
x"f6",
x"0d",
x"f2",
x"0b",
x"ce",
x"01",
x"03",
x"dd",
x"f2",
x"e1",
x"05",
x"03",
x"f7",
x"0e",
x"bb",
x"f7",
x"05",
x"e3",
x"fa",
x"e3",
x"f6",
x"f8",
x"f2",
x"06",
x"cd",
x"02",
x"fd",
x"f3",
x"e8",
x"ba",
x"ea",
x"0b",
x"00",
x"f6",
x"d6",
x"f4",
x"0d",
x"fc",
x"eb",
x"04",
x"ff",
x"05",
x"f0",
x"00",
x"e2",
x"04",
x"f6",
x"ff",
x"e6",
x"0c",
x"13",
x"da",
x"fc",
x"0b",
x"d1",
x"d9",
x"0d",
x"f7",
x"cb",
x"10",
x"fb",
x"e6",
x"f8",
x"f6",
x"b3",
x"ec",
x"26",
x"ff",
x"c8",
x"01",
x"07",
x"ed",
x"f9",
x"01",
x"b5",
x"eb",
x"11",
x"10",
x"aa",
x"fb",
x"0f",
x"fa",
x"fb",
x"ef",
x"8e",
x"e4",
x"f4",
x"0e",
x"bf",
x"e9",
x"fe",
x"fc",
x"fa",
x"13",
x"bd",
x"d7",
x"e9",
x"17",
x"a6",
x"e1",
x"07",
x"ef",
x"f5",
x"f7",
x"c2",
x"96",
x"f2",
x"2c",
x"d9",
x"e4",
x"4a",
x"ca",
x"d3",
x"14",
x"ee",
x"d6",
x"b2",
x"f7",
x"f5",
x"1b",
x"43",
x"e4",
x"19",
x"c3",
x"f9",
x"d8",
x"d2",
x"fb",
x"06",
x"23",
x"24",
x"f1",
x"e5",
x"e8",
x"f7",
x"01",
x"e9",
x"e7",
x"f8",
x"09",
x"fd",
x"f6",
x"03",
x"f9",
x"f7",
x"f8",
x"fc",
x"f9",
x"09",
x"f9",
x"06",
x"fc",
x"fa",
x"07",
x"00",
x"03",
x"09",
x"04",
x"05",
x"00",
x"fb",
x"06",
x"fa",
x"f8",
x"05",
x"ff",
x"07",
x"fc",
x"ff",
x"05",
x"f4",
x"13",
x"fe",
x"f9",
x"fa",
x"d9",
x"ea",
x"11",
x"e5",
x"cf",
x"c6",
x"db",
x"05",
x"11",
x"03",
x"17",
x"dd",
x"c6",
x"cd",
x"a8",
x"ba",
x"e6",
x"00",
x"1f",
x"ea",
x"17",
x"ac",
x"f9",
x"9a",
x"b1",
x"9d",
x"00",
x"df",
x"ea",
x"ef",
x"00",
x"a1",
x"11",
x"91",
x"bd",
x"c7",
x"0d",
x"d9",
x"04",
x"eb",
x"f1",
x"e3",
x"fa",
x"b1",
x"ae",
x"b0",
x"0b",
x"d8",
x"fe",
x"e4",
x"03",
x"d6",
x"f3",
x"a6",
x"c2",
x"8d",
x"25",
x"c9",
x"ef",
x"db",
x"08",
x"cc",
x"fb",
x"a9",
x"b0",
x"81",
x"1e",
x"dd",
x"ff",
x"d4",
x"13",
x"cc",
x"fb",
x"92",
x"75",
x"9b",
x"12",
x"de",
x"ff",
x"c8",
x"fa",
x"e1",
x"07",
x"b6",
x"75",
x"a1",
x"0f",
x"d8",
x"09",
x"f0",
x"1a",
x"e6",
x"fc",
x"96",
x"bb",
x"b9",
x"22",
x"c7",
x"04",
x"fd",
x"10",
x"db",
x"0a",
x"a8",
x"c3",
x"ce",
x"0b",
x"dc",
x"10",
x"a3",
x"02",
x"d8",
x"06",
x"96",
x"c0",
x"df",
x"0b",
x"d8",
x"02",
x"94",
x"0b",
x"e9",
x"01",
x"91",
x"95",
x"eb",
x"f7",
x"de",
x"06",
x"9f",
x"ff",
x"f7",
x"06",
x"8a",
x"71",
x"e0",
x"f6",
x"c7",
x"13",
x"93",
x"01",
x"f3",
x"07",
x"a3",
x"68",
x"ed",
x"db",
x"ce",
x"09",
x"90",
x"03",
x"ef",
x"1b",
x"85",
x"69",
x"cb",
x"eb",
x"d4",
x"07",
x"90",
x"06",
x"e5",
x"1e",
x"81",
x"94",
x"c6",
x"05",
x"b8",
x"fb",
x"aa",
x"fa",
x"ee",
x"20",
x"b7",
x"ae",
x"d9",
x"e9",
x"c6",
x"f6",
x"bb",
x"ef",
x"e4",
x"3f",
x"b2",
x"d0",
x"c9",
x"e2",
x"bc",
x"15",
x"cd",
x"03",
x"ba",
x"44",
x"ca",
x"e0",
x"ad",
x"fc",
x"df",
x"35",
x"ee",
x"05",
x"a5",
x"12",
x"b8",
x"f1",
x"ae",
x"d0",
x"f3",
x"34",
x"eb",
x"ef",
x"de",
x"15",
x"d0",
x"ee",
x"d5",
x"e4",
x"da",
x"32",
x"fa",
x"e5",
x"c8",
x"ef",
x"07",
x"f7",
x"1f",
x"fc",
x"ea",
x"f8",
x"03",
x"e9",
x"e8",
x"ff",
x"04",
x"05",
x"1d",
x"fe",
x"ef",
x"fb",
x"02",
x"ff",
x"e5",
x"e9",
x"f8",
x"fc",
x"00",
x"fd",
x"fb",
x"fe",
x"04",
x"04",
x"00",
x"f8",
x"fd",
x"f7",
x"f7",
x"0a",
x"0a",
x"06",
x"00",
x"08",
x"08",
x"fa",
x"01",
x"fa",
x"ff",
x"09",
x"04",
x"04",
x"08",
x"0a",
x"03",
x"f9",
x"0b",
x"03",
x"f7",
x"f9",
x"09",
x"01",
x"04",
x"fd",
x"f6",
x"ff",
x"ff",
x"f8",
x"fb",
x"ec",
x"df",
x"f8",
x"f8",
x"f5",
x"f2",
x"14",
x"f6",
x"df",
x"e0",
x"cd",
x"f0",
x"df",
x"f9",
x"ca",
x"e2",
x"41",
x"db",
x"db",
x"dc",
x"f2",
x"ec",
x"cc",
x"01",
x"d8",
x"b4",
x"21",
x"b3",
x"b6",
x"b3",
x"d5",
x"d8",
x"d2",
x"ff",
x"dd",
x"8f",
x"1f",
x"a8",
x"ac",
x"8e",
x"e9",
x"84",
x"af",
x"fb",
x"ef",
x"b3",
x"04",
x"8e",
x"a0",
x"93",
x"c7",
x"a5",
x"a8",
x"ef",
x"05",
x"b6",
x"0e",
x"82",
x"a0",
x"9d",
x"bd",
x"90",
x"d6",
x"f8",
x"05",
x"ac",
x"10",
x"7a",
x"b0",
x"7b",
x"c0",
x"a6",
x"d8",
x"ec",
x"08",
x"92",
x"06",
x"91",
x"9b",
x"95",
x"bc",
x"7b",
x"f6",
x"e7",
x"00",
x"b4",
x"00",
x"82",
x"78",
x"55",
x"a5",
x"93",
x"f3",
x"d8",
x"f5",
x"a5",
x"18",
x"85",
x"7f",
x"57",
x"aa",
x"76",
x"e4",
x"d3",
x"05",
x"a3",
x"04",
x"8a",
x"91",
x"57",
x"a8",
x"61",
x"ca",
x"ce",
x"fd",
x"b4",
x"27",
x"92",
x"c1",
x"75",
x"a9",
x"9d",
x"fb",
x"cf",
x"13",
x"3c",
x"06",
x"a2",
x"c0",
x"8b",
x"d3",
x"83",
x"ee",
x"db",
x"17",
x"5e",
x"19",
x"ae",
x"95",
x"a9",
x"d7",
x"87",
x"e2",
x"ca",
x"0f",
x"a7",
x"18",
x"b2",
x"c2",
x"97",
x"d9",
x"93",
x"e0",
x"c5",
x"1d",
x"b8",
x"20",
x"bf",
x"ca",
x"83",
x"fe",
x"9d",
x"e1",
x"e1",
x"16",
x"80",
x"16",
x"d9",
x"c8",
x"ab",
x"00",
x"96",
x"ff",
x"e6",
x"e2",
x"9f",
x"33",
x"c0",
x"ec",
x"b8",
x"fe",
x"94",
x"00",
x"ec",
x"0d",
x"d3",
x"12",
x"e0",
x"ed",
x"c8",
x"13",
x"bd",
x"0f",
x"e3",
x"21",
x"e1",
x"08",
x"dd",
x"e9",
x"e6",
x"d6",
x"d5",
x"00",
x"f8",
x"fb",
x"0f",
x"1c",
x"f5",
x"f6",
x"f5",
x"00",
x"f5",
x"e4",
x"02",
x"f1",
x"f3",
x"10",
x"f7",
x"fb",
x"f7",
x"fe",
x"01",
x"f8",
x"03",
x"08",
x"00",
x"f0",
x"0a",
x"f9",
x"f7",
x"09",
x"01",
x"00",
x"06",
x"03",
x"fa",
x"f7",
x"06",
x"ff",
x"08",
x"03",
x"03",
x"02",
x"ff",
x"fe",
x"03",
x"fb",
x"05",
x"08",
x"09",
x"fd",
x"02",
x"f8",
x"08",
x"f6",
x"06",
x"07",
x"0a",
x"01",
x"fb",
x"01",
x"05",
x"07",
x"fd",
x"ff",
x"fb",
x"07",
x"fa",
x"05",
x"04",
x"06",
x"fb",
x"fe",
x"fa",
x"04",
x"f8",
x"09",
x"fd",
x"f9",
x"09",
x"03",
x"fd",
x"fb",
x"fd",
x"07",
x"08",
x"f6",
x"f4",
x"ef",
x"07",
x"f8",
x"05",
x"05",
x"fa",
x"20",
x"fe",
x"ff",
x"f0",
x"f8",
x"02",
x"e2",
x"e5",
x"01",
x"fd",
x"0d",
x"f1",
x"dd",
x"de",
x"ef",
x"f3",
x"dc",
x"e4",
x"ee",
x"fd",
x"fd",
x"cf",
x"de",
x"cb",
x"e9",
x"de",
x"cf",
x"dc",
x"cf",
x"05",
x"f0",
x"b8",
x"09",
x"cf",
x"f9",
x"ec",
x"c1",
x"d1",
x"da",
x"03",
x"06",
x"b6",
x"00",
x"e4",
x"f2",
x"d4",
x"c4",
x"d6",
x"cc",
x"fa",
x"01",
x"c2",
x"ed",
x"c1",
x"cb",
x"bb",
x"a6",
x"c1",
x"f8",
x"f7",
x"21",
x"b4",
x"f8",
x"d3",
x"e4",
x"bd",
x"b6",
x"b1",
x"05",
x"f0",
x"07",
x"81",
x"ee",
x"bf",
x"d8",
x"b9",
x"b0",
x"ae",
x"f6",
x"fa",
x"02",
x"8e",
x"f1",
x"ca",
x"d7",
x"b3",
x"9f",
x"a3",
x"d5",
x"f5",
x"58",
x"87",
x"9a",
x"c4",
x"d5",
x"b4",
x"a6",
x"9c",
x"87",
x"df",
x"2a",
x"7f",
x"e8",
x"bf",
x"d6",
x"c0",
x"90",
x"c8",
x"88",
x"f0",
x"20",
x"c6",
x"d9",
x"d7",
x"dd",
x"c5",
x"9a",
x"c5",
x"9e",
x"ef",
x"23",
x"c4",
x"da",
x"d8",
x"e6",
x"b1",
x"99",
x"ce",
x"90",
x"fd",
x"5f",
x"ae",
x"bf",
x"e6",
x"da",
x"c1",
x"ac",
x"d1",
x"c4",
x"f3",
x"35",
x"c9",
x"e3",
x"da",
x"ed",
x"e1",
x"ca",
x"d1",
x"c8",
x"05",
x"2a",
x"da",
x"f2",
x"ee",
x"f6",
x"e5",
x"e4",
x"cb",
x"c8",
x"f2",
x"fc",
x"e1",
x"10",
x"e6",
x"f5",
x"cc",
x"ef",
x"d9",
x"e2",
x"e5",
x"35",
x"dd",
x"06",
x"e9",
x"fe",
x"dd",
x"ea",
x"d1",
x"e1",
x"f5",
x"20",
x"d3",
x"fb",
x"e7",
x"08",
x"ee",
x"ed",
x"ea",
x"e7",
x"00",
x"2b",
x"e7",
x"d7",
x"02",
x"07",
x"f8",
x"05",
x"fe",
x"01",
x"f8",
x"02",
x"07",
x"fa",
x"f7",
x"fe",
x"fe",
x"04",
x"f8",
x"01",
x"09",
x"f6",
x"05",
x"f6",
x"00",
x"fd",
x"f9",
x"00",
x"fc",
x"00",
x"ff",
x"fe",
x"fa",
x"0a",
x"fa",
x"08",
x"01",
x"09",
x"02",
x"0a",
x"06",
x"fe",
x"f8",
x"f5"
);

constant mem_ram_b1_init : mem8_t := (
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff"
);

constant mem_ram_b2_init : mem8_t := (
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff"
);

constant mem_ram_b3_init : mem8_t := (
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"ff",
x"ff",
x"ff",
x"00",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff"
);

end neorv32_dmem_image;
